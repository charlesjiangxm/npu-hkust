/*Copyright 2020-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

module aq_core(
  input   [2  :0]  biu_cp0_coreid,
  input            biu_cp0_me_int,
  input            biu_cp0_ms_int,
  input            biu_cp0_mt_int,
  input   [39 :0]  biu_cp0_rvba,
  input            biu_cp0_se_int,
  input            biu_cp0_ss_int,
  input            biu_cp0_st_int,
  input            biu_ifu_arready,
  input   [127:0]  biu_ifu_rdata,
  input            biu_ifu_rid,
  input            biu_ifu_rlast,
  input   [1  :0]  biu_ifu_rresp,
  input            biu_ifu_rvalid,
  input            biu_lsu_arready,
  input            biu_lsu_no_op,
  input   [127:0]  biu_lsu_rdata,
  input   [3  :0]  biu_lsu_rid,
  input            biu_lsu_rlast,
  input   [1  :0]  biu_lsu_rresp,
  input            biu_lsu_rvalid,
  input            biu_lsu_stb_awready,
  input            biu_lsu_stb_wready,
  input            biu_lsu_vb_awready,
  input            biu_lsu_vb_wready,
  input            cpurst_b,
  input            dtu_cp0_dcsr_mprven,
  input   [1  :0]  dtu_cp0_dcsr_prv,
  input   [63 :0]  dtu_cp0_rdata,
  input            dtu_cp0_wake_up,
  input   [31 :0]  dtu_ifu_debug_inst,
  input            dtu_ifu_debug_inst_vld,
  input   [21 :0]  dtu_ifu_halt_info0,
  input   [21 :0]  dtu_ifu_halt_info1,
  input            dtu_ifu_halt_info_vld,
  input            dtu_ifu_halt_on_reset,
  input            dtu_lsu_addr_trig_en,
  input            dtu_lsu_data_trig_en,
  input   [21 :0]  dtu_lsu_halt_info,
  input            dtu_lsu_halt_info_vld,
  input            dtu_rtu_async_halt_req,
  input   [63 :0]  dtu_rtu_dpc,
  input            dtu_rtu_ebreak_action,
  input            dtu_rtu_int_mask,
  input   [63 :0]  dtu_rtu_pending_tval,
  input            dtu_rtu_resume_req,
  input            dtu_rtu_step_en,
  input            dtu_rtu_sync_flush,
  input            dtu_rtu_sync_halt_req,
  input            forever_cpuclk,
  input   [63 :0]  hpcp_cp0_data,
  input            hpcp_cp0_int_vld,
  input            hpcp_cp0_sce,
  input            hpcp_idu_cnt_en,
  input            hpcp_ifu_cnt_en,
  input            hpcp_iu_cnt_en,
  input            hpcp_lsu_cnt_en,
  input            hpcp_rtu_cnt_en,
  input            mmu_cp0_cmplt,
  input   [63 :0]  mmu_cp0_data,
  input            mmu_cp0_tlb_inv_done,
  input            mmu_ifu_access_fault,
  input   [27 :0]  mmu_ifu_pa,
  input            mmu_ifu_pa_vld,
  input   [4  :0]  mmu_ifu_prot,
  input            mmu_lsu_access_fault,
  input            mmu_lsu_buf,
  input            mmu_lsu_ca,
  input            mmu_lsu_data_req,
  input   [39 :0]  mmu_lsu_data_req_addr,
  input            mmu_lsu_data_req_size,
  input   [27 :0]  mmu_lsu_pa,
  input            mmu_lsu_pa_vld,
  input            mmu_lsu_page_fault,
  input            mmu_lsu_sec,
  input            mmu_lsu_sh,
  input            mmu_lsu_so,
  input            mmu_xx_mmu_en,
  input            mmu_yy_xx_no_op,
  input            pad_yy_icg_scan_en,
  input            pad_yy_scan_mode,
  input   [63 :0]  pmp_cp0_data,
  input   [39 :0]  sysio_cp0_apb_base,
  output           cp0_biu_icg_en,
  output  [1  :0]  cp0_biu_lpmd_b,
  output  [11 :0]  cp0_dtu_addr,
  output  [5  :0]  cp0_dtu_debug_info,
  output           cp0_dtu_icg_en,
  output           cp0_dtu_mexpt_vld,
  output           cp0_dtu_pcfifo_frz,
  output           cp0_dtu_rreg,
  output  [63 :0]  cp0_dtu_satp,
  output  [63 :0]  cp0_dtu_wdata,
  output           cp0_dtu_wreg,
  output           cp0_hpcp_icg_en,
  output  [11 :0]  cp0_hpcp_index,
  output           cp0_hpcp_int_off_vld,
  output  [31 :0]  cp0_hpcp_mcntwen,
  output           cp0_hpcp_pmdm,
  output           cp0_hpcp_pmds,
  output           cp0_hpcp_pmdu,
  output           cp0_hpcp_sync_stall_vld,
  output  [63 :0]  cp0_hpcp_wdata,
  output           cp0_hpcp_wreg,
  output  [11 :0]  cp0_mmu_addr,
  output           cp0_mmu_icg_en,
  output           cp0_mmu_lpmd_req,
  output           cp0_mmu_maee,
  output           cp0_mmu_mxr,
  output           cp0_mmu_ptw_en,
  output  [63 :0]  cp0_mmu_satp_data,
  output           cp0_mmu_satp_wen,
  output           cp0_mmu_sum,
  output           cp0_mmu_tlb_all_inv,
  output  [15 :0]  cp0_mmu_tlb_asid,
  output           cp0_mmu_tlb_asid_all_inv,
  output  [26 :0]  cp0_mmu_tlb_va,
  output           cp0_mmu_tlb_va_all_inv,
  output           cp0_mmu_tlb_va_asid_inv,
  output  [63 :0]  cp0_mmu_wdata,
  output           cp0_mmu_wreg,
  output  [11 :0]  cp0_pmp_addr,
  output           cp0_pmp_icg_en,
  output  [63 :0]  cp0_pmp_wdata,
  output           cp0_pmp_wreg,
  output           cp0_yy_clk_en,
  output  [1  :0]  cp0_yy_priv_mode,
  output  [14 :0]  idu_dtu_debug_info,
  output           idu_hpcp_backend_stall,
  output           idu_hpcp_frontend_stall,
  output  [6  :0]  idu_hpcp_inst_type,
  output  [39 :0]  ifu_biu_araddr,
  output  [1  :0]  ifu_biu_arburst,
  output  [3  :0]  ifu_biu_arcache,
  output           ifu_biu_arid,
  output  [1  :0]  ifu_biu_arlen,
  output  [2  :0]  ifu_biu_arprot,
  output  [2  :0]  ifu_biu_arsize,
  output           ifu_biu_arvalid,
  output           ifu_dtu_addr_vld0,
  output           ifu_dtu_addr_vld1,
  output           ifu_dtu_data_vld0,
  output           ifu_dtu_data_vld1,
  output  [20 :0]  ifu_dtu_debug_info,
  output  [39 :0]  ifu_dtu_exe_addr0,
  output  [39 :0]  ifu_dtu_exe_addr1,
  output  [31 :0]  ifu_dtu_exe_data0,
  output  [31 :0]  ifu_dtu_exe_data1,
  output           ifu_hpcp_icache_access,
  output           ifu_hpcp_icache_miss,
  output           ifu_mmu_abort,
  output  [51 :0]  ifu_mmu_va,
  output           ifu_mmu_va_vld,
  output  [8  :0]  iu_dtu_debug_info,
  output           iu_hpcp_inst_bht_mispred,
  output           iu_hpcp_inst_condbr,
  output           iu_hpcp_jump_8m,
  output  [39 :0]  lsu_biu_araddr,
  output  [1  :0]  lsu_biu_arburst,
  output  [3  :0]  lsu_biu_arcache,
  output  [3  :0]  lsu_biu_arid,
  output  [1  :0]  lsu_biu_arlen,
  output  [2  :0]  lsu_biu_arprot,
  output  [2  :0]  lsu_biu_arsize,
  output           lsu_biu_aruser,
  output           lsu_biu_arvalid,
  output  [39 :0]  lsu_biu_stb_awaddr,
  output  [1  :0]  lsu_biu_stb_awburst,
  output  [3  :0]  lsu_biu_stb_awcache,
  output  [1  :0]  lsu_biu_stb_awid,
  output  [1  :0]  lsu_biu_stb_awlen,
  output  [2  :0]  lsu_biu_stb_awprot,
  output  [2  :0]  lsu_biu_stb_awsize,
  output           lsu_biu_stb_awuser,
  output           lsu_biu_stb_awvalid,
  output  [127:0]  lsu_biu_stb_wdata,
  output           lsu_biu_stb_wlast,
  output  [15 :0]  lsu_biu_stb_wstrb,
  output           lsu_biu_stb_wvalid,
  output  [39 :0]  lsu_biu_vb_awaddr,
  output  [1  :0]  lsu_biu_vb_awburst,
  output  [3  :0]  lsu_biu_vb_awcache,
  output  [3  :0]  lsu_biu_vb_awid,
  output  [1  :0]  lsu_biu_vb_awlen,
  output  [2  :0]  lsu_biu_vb_awprot,
  output  [2  :0]  lsu_biu_vb_awsize,
  output           lsu_biu_vb_awvalid,
  output  [127:0]  lsu_biu_vb_wdata,
  output           lsu_biu_vb_wlast,
  output  [15 :0]  lsu_biu_vb_wstrb,
  output           lsu_biu_vb_wvalid,
  output  [93 :0]  lsu_dtu_debug_info,
  output  [21 :0]  lsu_dtu_halt_info,
  output           lsu_dtu_last_check,
  output  [39 :0]  lsu_dtu_ldst_addr,
  output           lsu_dtu_ldst_addr_vld,
  output  [15 :0]  lsu_dtu_ldst_bytes_vld,
  output  [63 :0]  lsu_dtu_ldst_data,
  output           lsu_dtu_ldst_data_vld,
  output  [1  :0]  lsu_dtu_ldst_type,
  output  [2  :0]  lsu_dtu_mem_access_size,
  output           lsu_hpcp_cache_read_access,
  output           lsu_hpcp_cache_read_miss,
  output           lsu_hpcp_cache_write_access,
  output           lsu_hpcp_cache_write_miss,
  output           lsu_hpcp_inst_store,
  output           lsu_hpcp_unalign_inst,
  output           lsu_mmu_abort,
  output           lsu_mmu_bus_error,
  output  [63 :0]  lsu_mmu_data,
  output           lsu_mmu_data_vld,
  output  [1  :0]  lsu_mmu_priv_mode,
  output           lsu_mmu_st_inst,
  output  [51 :0]  lsu_mmu_va,
  output           lsu_mmu_va_vld,
  output           rtu_cpu_no_retire,
  output  [14 :0]  rtu_dtu_debug_info,
  output  [63 :0]  rtu_dtu_dpc,
  output           rtu_dtu_halt_ack,
  output           rtu_dtu_pending_ack,
  output           rtu_dtu_retire_chgflw,
  output           rtu_dtu_retire_debug_expt_vld,
  output  [21 :0]  rtu_dtu_retire_halt_info,
  output           rtu_dtu_retire_mret,
  output  [39 :0]  rtu_dtu_retire_next_pc,
  output           rtu_dtu_retire_sret,
  output           rtu_dtu_retire_vld,
  output  [63 :0]  rtu_dtu_tval,
  output           rtu_hpcp_int_vld,
  output           rtu_hpcp_retire_inst_vld,
  output  [39 :0]  rtu_hpcp_retire_pc,
  output  [26 :0]  rtu_mmu_bad_vpn,
  output           rtu_mmu_expt_vld,
  output           rtu_pad_halted,
  output           rtu_pad_retire,
  output  [39 :0]  rtu_pad_retire_pc,
  output           rtu_yy_xx_dbgon,
  output           rtu_yy_xx_expt_int,
  output  [4  :0]  rtu_yy_xx_expt_vec,
  output           rtu_yy_xx_expt_vld,
  output  [7  :0]  vidu_dtu_debug_info,
  output  [28 :0]  vpu_dtu_dbg_info
);

aq_ifu_top  x_aq_ifu_top (
  .biu_ifu_arready              (biu_ifu_arready             ),
  .biu_ifu_rdata                (biu_ifu_rdata               ),
  .biu_ifu_rid                  (biu_ifu_rid                 ),
  .biu_ifu_rlast                (biu_ifu_rlast               ),
  .biu_ifu_rresp                (biu_ifu_rresp               ),
  .biu_ifu_rvalid               (biu_ifu_rvalid              ),
  .cp0_ifu_bht_en               (cp0_ifu_bht_en              ),
  .cp0_ifu_bht_inv              (cp0_ifu_bht_inv             ),
  .cp0_ifu_btb_clr              (cp0_ifu_btb_clr             ),
  .cp0_ifu_btb_en               (cp0_ifu_btb_en              ),
  .cp0_ifu_icache_en            (cp0_ifu_icache_en           ),
  .cp0_ifu_icache_inv_addr      (cp0_ifu_icache_inv_addr     ),
  .cp0_ifu_icache_inv_req       (cp0_ifu_icache_inv_req      ),
  .cp0_ifu_icache_inv_type      (cp0_ifu_icache_inv_type     ),
  .cp0_ifu_icache_pref_en       (cp0_ifu_icache_pref_en      ),
  .cp0_ifu_icache_read_index    (cp0_ifu_icache_read_index   ),
  .cp0_ifu_icache_read_req      (cp0_ifu_icache_read_req     ),
  .cp0_ifu_icache_read_tag      (cp0_ifu_icache_read_tag     ),
  .cp0_ifu_icache_read_way      (cp0_ifu_icache_read_way     ),
  .cp0_ifu_icg_en               (cp0_ifu_icg_en              ),
  .cp0_ifu_in_lpmd              (cp0_ifu_in_lpmd             ),
  .cp0_ifu_iwpe                 (cp0_ifu_iwpe                ),
  .cp0_ifu_lpmd_req             (cp0_ifu_lpmd_req            ),
  .cp0_ifu_ras_en               (cp0_ifu_ras_en              ),
  .cp0_ifu_rst_inv_done         (cp0_ifu_rst_inv_done        ),
  .cp0_xx_mrvbr                 (cp0_xx_mrvbr                ),
  .cp0_yy_clk_en                (cp0_yy_clk_en               ),
  .cpurst_b                     (cpurst_b                    ),
  .dtu_ifu_debug_inst           (dtu_ifu_debug_inst          ),
  .dtu_ifu_debug_inst_vld       (dtu_ifu_debug_inst_vld      ),
  .dtu_ifu_halt_info0           (dtu_ifu_halt_info0          ),
  .dtu_ifu_halt_info1           (dtu_ifu_halt_info1          ),
  .dtu_ifu_halt_info_vld        (dtu_ifu_halt_info_vld       ),
  .dtu_ifu_halt_on_reset        (dtu_ifu_halt_on_reset       ),
  .forever_cpuclk               (forever_cpuclk              ),
  .hpcp_ifu_cnt_en              (hpcp_ifu_cnt_en             ),
  .idu_ifu_id_stall             (idu_ifu_id_stall            ),
  .ifu_biu_araddr               (ifu_biu_araddr              ),
  .ifu_biu_arburst              (ifu_biu_arburst             ),
  .ifu_biu_arcache              (ifu_biu_arcache             ),
  .ifu_biu_arid                 (ifu_biu_arid                ),
  .ifu_biu_arlen                (ifu_biu_arlen               ),
  .ifu_biu_arprot               (ifu_biu_arprot              ),
  .ifu_biu_arsize               (ifu_biu_arsize              ),
  .ifu_biu_arvalid              (ifu_biu_arvalid             ),
  .ifu_cp0_bht_inv_done         (ifu_cp0_bht_inv_done        ),
  .ifu_cp0_icache_inv_done      (ifu_cp0_icache_inv_done     ),
  .ifu_cp0_icache_read_data     (ifu_cp0_icache_read_data    ),
  .ifu_cp0_icache_read_data_vld (ifu_cp0_icache_read_data_vld),
  .ifu_cp0_rst_inv_req          (ifu_cp0_rst_inv_req         ),
  .ifu_cp0_warm_up              (ifu_cp0_warm_up             ),
  .ifu_dtu_addr_vld0            (ifu_dtu_addr_vld0           ),
  .ifu_dtu_addr_vld1            (ifu_dtu_addr_vld1           ),
  .ifu_dtu_data_vld0            (ifu_dtu_data_vld0           ),
  .ifu_dtu_data_vld1            (ifu_dtu_data_vld1           ),
  .ifu_dtu_debug_info           (ifu_dtu_debug_info          ),
  .ifu_dtu_exe_addr0            (ifu_dtu_exe_addr0           ),
  .ifu_dtu_exe_addr1            (ifu_dtu_exe_addr1           ),
  .ifu_dtu_exe_data0            (ifu_dtu_exe_data0           ),
  .ifu_dtu_exe_data1            (ifu_dtu_exe_data1           ),
  .ifu_hpcp_icache_access       (ifu_hpcp_icache_access      ),
  .ifu_hpcp_icache_miss         (ifu_hpcp_icache_miss        ),
  .ifu_idu_id_bht_pred          (ifu_idu_id_bht_pred         ),
  .ifu_idu_id_expt_acc_error    (ifu_idu_id_expt_acc_error   ),
  .ifu_idu_id_expt_high         (ifu_idu_id_expt_high        ),
  .ifu_idu_id_expt_page_fault   (ifu_idu_id_expt_page_fault  ),
  .ifu_idu_id_halt_info         (ifu_idu_id_halt_info        ),
  .ifu_idu_id_inst              (ifu_idu_id_inst             ),
  .ifu_idu_id_inst_vld          (ifu_idu_id_inst_vld         ),
  .ifu_idu_warm_up              (ifu_idu_warm_up             ),
  .ifu_iu_chgflw_pc             (ifu_iu_chgflw_pc            ),
  .ifu_iu_chgflw_vld            (ifu_iu_chgflw_vld           ),
  .ifu_iu_ex1_pc_pred           (ifu_iu_ex1_pc_pred          ),
  .ifu_iu_reset_vld             (ifu_iu_reset_vld            ),
  .ifu_iu_warm_up               (ifu_iu_warm_up              ),
  .ifu_lsu_warm_up              (ifu_lsu_warm_up             ),
  .ifu_mmu_abort                (ifu_mmu_abort               ),
  .ifu_mmu_va                   (ifu_mmu_va                  ),
  .ifu_mmu_va_vld               (ifu_mmu_va_vld              ),
  .ifu_rtu_reset_halt_req       (ifu_rtu_reset_halt_req      ),
  .ifu_rtu_warm_up              (ifu_rtu_warm_up             ),
  .ifu_vidu_warm_up             (ifu_vidu_warm_up            ),
  .ifu_vpu_warm_up              (ifu_vpu_warm_up             ),
  .ifu_yy_xx_no_op              (ifu_yy_xx_no_op             ),
  .iu_ifu_bht_cur_pc            (iu_ifu_bht_cur_pc           ),
  .iu_ifu_bht_mispred           (iu_ifu_bht_mispred          ),
  .iu_ifu_bht_mispred_gate      (iu_ifu_bht_mispred_gate     ),
  .iu_ifu_bht_pred              (iu_ifu_bht_pred             ),
  .iu_ifu_bht_taken             (iu_ifu_bht_taken            ),
  .iu_ifu_br_vld                (iu_ifu_br_vld               ),
  .iu_ifu_br_vld_gate           (iu_ifu_br_vld_gate          ),
  .iu_ifu_link_vld              (iu_ifu_link_vld             ),
  .iu_ifu_link_vld_gate         (iu_ifu_link_vld_gate        ),
  .iu_ifu_pc_mispred            (iu_ifu_pc_mispred           ),
  .iu_ifu_pc_mispred_gate       (iu_ifu_pc_mispred_gate      ),
  .iu_ifu_ret_vld               (iu_ifu_ret_vld              ),
  .iu_ifu_ret_vld_gate          (iu_ifu_ret_vld_gate         ),
  .iu_ifu_tar_pc                (iu_ifu_tar_pc               ),
  .iu_ifu_tar_pc_vld            (iu_ifu_tar_pc_vld           ),
  .iu_ifu_tar_pc_vld_gate       (iu_ifu_tar_pc_vld_gate      ),
  .mmu_ifu_access_fault         (mmu_ifu_access_fault        ),
  .mmu_ifu_pa                   (mmu_ifu_pa                  ),
  .mmu_ifu_pa_vld               (mmu_ifu_pa_vld              ),
  .mmu_ifu_prot                 (mmu_ifu_prot                ),
  .pad_yy_icg_scan_en           (pad_yy_icg_scan_en          ),
  .rtu_ifu_chgflw_pc            (rtu_ifu_chgflw_pc           ),
  .rtu_ifu_chgflw_vld           (rtu_ifu_chgflw_vld          ),
  .rtu_ifu_dbg_mask             (rtu_ifu_dbg_mask            ),
  .rtu_ifu_flush_fe             (rtu_ifu_flush_fe            ),
  .rtu_yy_xx_dbgon              (rtu_yy_xx_dbgon             )
);


aq_idu_top  x_aq_idu_top (
  .cp0_idu_cskyee               (cp0_idu_cskyee              ),
  .cp0_idu_dis_fence_in_dbg     (cp0_idu_dis_fence_in_dbg    ),
  .cp0_idu_frm                  (cp0_idu_frm                 ),
  .cp0_idu_fs                   (cp0_idu_fs                  ),
  .cp0_idu_icg_en               (cp0_idu_icg_en              ),
  .cp0_idu_issue_stall          (cp0_idu_issue_stall         ),
  .cp0_idu_ucme                 (cp0_idu_ucme                ),
  .cp0_idu_vill                 (cp0_idu_vill                ),
  .cp0_idu_vl_zero              (cp0_idu_vl_zero             ),
  .cp0_idu_vlmul                (cp0_idu_vlmul               ),
  .cp0_idu_vs                   (cp0_idu_vs                  ),
  .cp0_idu_vsetvl_dis_stall     (cp0_idu_vsetvl_dis_stall    ),
  .cp0_idu_vsew                 (cp0_idu_vsew                ),
  .cp0_idu_vstart               (cp0_idu_vstart              ),
  .cp0_yy_clk_en                (cp0_yy_clk_en               ),
  .cp0_yy_priv_mode             (cp0_yy_priv_mode            ),
  .cpurst_b                     (cpurst_b                    ),
  .forever_cpuclk               (forever_cpuclk              ),
  .hpcp_idu_cnt_en              (hpcp_idu_cnt_en             ),
  .idu_alu_ex1_gateclk_sel      (idu_alu_ex1_gateclk_sel     ),
  .idu_bju_ex1_gateclk_sel      (idu_bju_ex1_gateclk_sel     ),
  .idu_cp0_ex1_dp_sel           (idu_cp0_ex1_dp_sel          ),
  .idu_cp0_ex1_dst0_reg         (idu_cp0_ex1_dst0_reg        ),
  .idu_cp0_ex1_expt_acc_error   (idu_cp0_ex1_expt_acc_error  ),
  .idu_cp0_ex1_expt_high        (idu_cp0_ex1_expt_high       ),
  .idu_cp0_ex1_expt_illegal     (idu_cp0_ex1_expt_illegal    ),
  .idu_cp0_ex1_expt_page_fault  (idu_cp0_ex1_expt_page_fault ),
  .idu_cp0_ex1_func             (idu_cp0_ex1_func            ),
  .idu_cp0_ex1_gateclk_sel      (idu_cp0_ex1_gateclk_sel     ),
  .idu_cp0_ex1_halt_info        (idu_cp0_ex1_halt_info       ),
  .idu_cp0_ex1_length           (idu_cp0_ex1_length          ),
  .idu_cp0_ex1_opcode           (idu_cp0_ex1_opcode          ),
  .idu_cp0_ex1_sel              (idu_cp0_ex1_sel             ),
  .idu_cp0_ex1_split            (idu_cp0_ex1_split           ),
  .idu_cp0_ex1_src0_data        (idu_cp0_ex1_src0_data       ),
  .idu_cp0_ex1_src1_data        (idu_cp0_ex1_src1_data       ),
  .idu_div_ex1_gateclk_sel      (idu_div_ex1_gateclk_sel     ),
  .idu_dtu_debug_info           (idu_dtu_debug_info          ),
  .idu_hpcp_backend_stall       (idu_hpcp_backend_stall      ),
  .idu_hpcp_frontend_stall      (idu_hpcp_frontend_stall     ),
  .idu_hpcp_inst_type           (idu_hpcp_inst_type          ),
  .idu_ifu_id_stall             (idu_ifu_id_stall            ),
  .idu_iu_ex1_alu_dp_sel        (idu_iu_ex1_alu_dp_sel       ),
  .idu_iu_ex1_alu_sel           (idu_iu_ex1_alu_sel          ),
  .idu_iu_ex1_bht_pred          (idu_iu_ex1_bht_pred         ),
  .idu_iu_ex1_bju_br_sel        (idu_iu_ex1_bju_br_sel       ),
  .idu_iu_ex1_bju_dp_sel        (idu_iu_ex1_bju_dp_sel       ),
  .idu_iu_ex1_bju_sel           (idu_iu_ex1_bju_sel          ),
  .idu_iu_ex1_div_dp_sel        (idu_iu_ex1_div_dp_sel       ),
  .idu_iu_ex1_div_sel           (idu_iu_ex1_div_sel          ),
  .idu_iu_ex1_dst0_reg          (idu_iu_ex1_dst0_reg         ),
  .idu_iu_ex1_func              (idu_iu_ex1_func             ),
  .idu_iu_ex1_inst_vld          (idu_iu_ex1_inst_vld         ),
  .idu_iu_ex1_length            (idu_iu_ex1_length           ),
  .idu_iu_ex1_mult_dp_sel       (idu_iu_ex1_mult_dp_sel      ),
  .idu_iu_ex1_mult_sel          (idu_iu_ex1_mult_sel         ),
  .idu_iu_ex1_pipedown_vld      (idu_iu_ex1_pipedown_vld     ),
  .idu_iu_ex1_split             (idu_iu_ex1_split            ),
  .idu_iu_ex1_src0_data         (idu_iu_ex1_src0_data        ),
  .idu_iu_ex1_src0_ready        (idu_iu_ex1_src0_ready       ),
  .idu_iu_ex1_src0_reg          (idu_iu_ex1_src0_reg         ),
  .idu_iu_ex1_src1_data         (idu_iu_ex1_src1_data        ),
  .idu_iu_ex1_src1_ready        (idu_iu_ex1_src1_ready       ),
  .idu_iu_ex1_src1_reg          (idu_iu_ex1_src1_reg         ),
  .idu_iu_ex1_src2_data         (idu_iu_ex1_src2_data        ),
  .idu_lsu_ex1_dp_sel           (idu_lsu_ex1_dp_sel          ),
  .idu_lsu_ex1_dst0_reg         (idu_lsu_ex1_dst0_reg        ),
  .idu_lsu_ex1_dst1_reg         (idu_lsu_ex1_dst1_reg        ),
  .idu_lsu_ex1_func             (idu_lsu_ex1_func            ),
  .idu_lsu_ex1_gateclk_sel      (idu_lsu_ex1_gateclk_sel     ),
  .idu_lsu_ex1_halt_info        (idu_lsu_ex1_halt_info       ),
  .idu_lsu_ex1_length           (idu_lsu_ex1_length          ),
  .idu_lsu_ex1_sel              (idu_lsu_ex1_sel             ),
  .idu_lsu_ex1_split            (idu_lsu_ex1_split           ),
  .idu_lsu_ex1_src0_data        (idu_lsu_ex1_src0_data       ),
  .idu_lsu_ex1_src1_data        (idu_lsu_ex1_src1_data       ),
  .idu_lsu_ex1_src2_data        (idu_lsu_ex1_src2_data       ),
  .idu_lsu_ex1_src2_ready       (idu_lsu_ex1_src2_ready      ),
  .idu_lsu_ex1_src2_reg         (idu_lsu_ex1_src2_reg        ),
  .idu_lsu_ex1_vlmul            (idu_lsu_ex1_vlmul           ),
  .idu_lsu_ex1_vsew             (idu_lsu_ex1_vsew            ),
  .idu_mult_ex1_gateclk_sel     (idu_mult_ex1_gateclk_sel    ),
  .idu_vidu_ex1_fp_dp_sel       (idu_vidu_ex1_fp_dp_sel      ),
  .idu_vidu_ex1_fp_gateclk_sel  (idu_vidu_ex1_fp_gateclk_sel ),
  .idu_vidu_ex1_fp_sel          (idu_vidu_ex1_fp_sel         ),
  .idu_vidu_ex1_inst_data       (idu_vidu_ex1_inst_data      ),
  .idu_vidu_ex1_vec_dp_sel      (idu_vidu_ex1_vec_dp_sel     ),
  .idu_vidu_ex1_vec_gateclk_sel (idu_vidu_ex1_vec_gateclk_sel),
  .idu_vidu_ex1_vec_sel         (idu_vidu_ex1_vec_sel        ),
  .ifu_idu_id_bht_pred          (ifu_idu_id_bht_pred         ),
  .ifu_idu_id_expt_acc_error    (ifu_idu_id_expt_acc_error   ),
  .ifu_idu_id_expt_high         (ifu_idu_id_expt_high        ),
  .ifu_idu_id_expt_page_fault   (ifu_idu_id_expt_page_fault  ),
  .ifu_idu_id_halt_info         (ifu_idu_id_halt_info        ),
  .ifu_idu_id_inst              (ifu_idu_id_inst             ),
  .ifu_idu_id_inst_vld          (ifu_idu_id_inst_vld         ),
  .ifu_idu_warm_up              (ifu_idu_warm_up             ),
  .iu_idu_bju_full              (iu_idu_bju_full             ),
  .iu_idu_bju_global_full       (iu_idu_bju_global_full      ),
  .iu_idu_div_full              (iu_idu_div_full             ),
  .iu_idu_mult_full             (iu_idu_mult_full            ),
  .iu_idu_mult_issue_stall      (iu_idu_mult_issue_stall     ),
  .iu_yy_xx_cancel              (iu_yy_xx_cancel             ),
  .lsu_idu_full                 (lsu_idu_full                ),
  .lsu_idu_global_full          (lsu_idu_global_full         ),
  .pad_yy_icg_scan_en           (pad_yy_icg_scan_en          ),
  .rtu_idu_commit               (rtu_idu_commit              ),
  .rtu_idu_commit_for_bju       (rtu_idu_commit_for_bju      ),
  .rtu_idu_flush_fe             (rtu_idu_flush_fe            ),
  .rtu_idu_flush_stall          (rtu_idu_flush_stall         ),
  .rtu_idu_flush_wbt            (rtu_idu_flush_wbt           ),
  .rtu_idu_fwd0_data            (rtu_idu_fwd0_data           ),
  .rtu_idu_fwd0_reg             (rtu_idu_fwd0_reg            ),
  .rtu_idu_fwd0_vld             (rtu_idu_fwd0_vld            ),
  .rtu_idu_fwd1_data            (rtu_idu_fwd1_data           ),
  .rtu_idu_fwd1_reg             (rtu_idu_fwd1_reg            ),
  .rtu_idu_fwd1_vld             (rtu_idu_fwd1_vld            ),
  .rtu_idu_fwd2_data            (rtu_idu_fwd2_data           ),
  .rtu_idu_fwd2_reg             (rtu_idu_fwd2_reg            ),
  .rtu_idu_fwd2_vld             (rtu_idu_fwd2_vld            ),
  .rtu_idu_pipeline_empty       (rtu_idu_pipeline_empty      ),
  .rtu_idu_wb0_data             (rtu_idu_wb0_data            ),
  .rtu_idu_wb0_reg              (rtu_idu_wb0_reg             ),
  .rtu_idu_wb0_vld              (rtu_idu_wb0_vld             ),
  .rtu_idu_wb1_data             (rtu_idu_wb1_data            ),
  .rtu_idu_wb1_reg              (rtu_idu_wb1_reg             ),
  .rtu_idu_wb1_vld              (rtu_idu_wb1_vld             ),
  .rtu_yy_xx_dbgon              (rtu_yy_xx_dbgon             ),
  .vidu_idu_fp_full             (vidu_idu_fp_full            ),
  .vidu_idu_vec_full            (vidu_idu_vec_full           )
);

aq_vidu_top  x_aq_vidu_top (
  .cp0_idu_icg_en                   (cp0_idu_icg_en                  ),
  .cp0_yy_clk_en                    (cp0_yy_clk_en                   ),
  .cpurst_b                         (cpurst_b                        ),
  .forever_cpuclk                   (forever_cpuclk                  ),
  .idu_vidu_ex1_fp_dp_sel           (idu_vidu_ex1_fp_dp_sel          ),
  .idu_vidu_ex1_fp_gateclk_sel      (idu_vidu_ex1_fp_gateclk_sel     ),
  .idu_vidu_ex1_fp_sel              (idu_vidu_ex1_fp_sel             ),
  .idu_vidu_ex1_inst_data           (idu_vidu_ex1_inst_data          ),
  .idu_vidu_ex1_vec_dp_sel          (idu_vidu_ex1_vec_dp_sel         ),
  .idu_vidu_ex1_vec_gateclk_sel     (idu_vidu_ex1_vec_gateclk_sel    ),
  .idu_vidu_ex1_vec_sel             (idu_vidu_ex1_vec_sel            ),
  .ifu_vidu_warm_up                 (ifu_vidu_warm_up                ),
  .pad_yy_icg_scan_en               (pad_yy_icg_scan_en              ),
  .rtu_vidu_flush_wbt               (rtu_vidu_flush_wbt              ),
  .rtu_yy_xx_async_flush            (rtu_yy_xx_async_flush           ),
  .vidu_cp0_vid_fof_vld             (vidu_cp0_vid_fof_vld            ),
  .vidu_dtu_debug_info              (vidu_dtu_debug_info             ),
  .vidu_idu_fp_full                 (vidu_idu_fp_full                ),
  .vidu_idu_vec_full                (vidu_idu_vec_full               ),
  .vidu_rtu_no_op                   (vidu_rtu_no_op                  ),
  .vidu_vpu_vid_fp_inst_dp_vld      (vidu_vpu_vid_fp_inst_dp_vld     ),
  .vidu_vpu_vid_fp_inst_dst_reg     (vidu_vpu_vid_fp_inst_dst_reg    ),
  .vidu_vpu_vid_fp_inst_dst_vld     (vidu_vpu_vid_fp_inst_dst_vld    ),
  .vidu_vpu_vid_fp_inst_dste_vld    (vidu_vpu_vid_fp_inst_dste_vld   ),
  .vidu_vpu_vid_fp_inst_dstf_reg    (vidu_vpu_vid_fp_inst_dstf_reg   ),
  .vidu_vpu_vid_fp_inst_dstf_vld    (vidu_vpu_vid_fp_inst_dstf_vld   ),
  .vidu_vpu_vid_fp_inst_eu          (vidu_vpu_vid_fp_inst_eu         ),
  .vidu_vpu_vid_fp_inst_func        (vidu_vpu_vid_fp_inst_func       ),
  .vidu_vpu_vid_fp_inst_gateclk_vld (vidu_vpu_vid_fp_inst_gateclk_vld),
  .vidu_vpu_vid_fp_inst_src1_data   (vidu_vpu_vid_fp_inst_src1_data  ),
  .vidu_vpu_vid_fp_inst_srcf0_data  (vidu_vpu_vid_fp_inst_srcf0_data ),
  .vidu_vpu_vid_fp_inst_srcf1_data  (vidu_vpu_vid_fp_inst_srcf1_data ),
  .vidu_vpu_vid_fp_inst_srcf2_data  (vidu_vpu_vid_fp_inst_srcf2_data ),
  .vidu_vpu_vid_fp_inst_srcf2_rdy   (vidu_vpu_vid_fp_inst_srcf2_rdy  ),
  .vidu_vpu_vid_fp_inst_srcf2_vld   (vidu_vpu_vid_fp_inst_srcf2_vld  ),
  .vidu_vpu_vid_fp_inst_vld         (vidu_vpu_vid_fp_inst_vld        ),
  .vpu_rtu_ex1_cmplt                (vpu_rtu_ex1_cmplt               ),
  .vpu_rtu_ex1_cmplt_dp             (vpu_rtu_ex1_cmplt_dp            ),
  .vpu_rtu_ex1_fp_dirty             (vpu_rtu_ex1_fp_dirty            ),
  .vpu_rtu_ex1_vec_dirty            (vpu_rtu_ex1_vec_dirty           ),
  .vpu_vidu_fp_fwd_data             (vpu_vidu_fp_fwd_data            ),
  .vpu_vidu_fp_fwd_reg              (vpu_vidu_fp_fwd_reg             ),
  .vpu_vidu_fp_fwd_vld              (vpu_vidu_fp_fwd_vld             ),
  .vpu_vidu_fp_wb_data              (vpu_vidu_fp_wb_data             ),
  .vpu_vidu_fp_wb_reg               (vpu_vidu_fp_wb_reg              ),
  .vpu_vidu_fp_wb_vld               (vpu_vidu_fp_wb_vld              ),
  .vpu_vidu_vex1_fp_stall           (vpu_vidu_vex1_fp_stall          ),
  .vpu_vidu_wbt_fp_wb0_reg          (vpu_vidu_wbt_fp_wb0_reg         ),
  .vpu_vidu_wbt_fp_wb0_vld          (vpu_vidu_wbt_fp_wb0_vld         ),
  .vpu_vidu_wbt_fp_wb1_reg          (vpu_vidu_wbt_fp_wb1_reg         ),
  .vpu_vidu_wbt_fp_wb1_vld          (vpu_vidu_wbt_fp_wb1_vld         )
);

aq_iu_top  x_aq_iu_top (
  .cp0_iu_icg_en                (cp0_iu_icg_en               ),
  .cp0_xx_mrvbr                 (cp0_xx_mrvbr                ),
  .cp0_yy_clk_en                (cp0_yy_clk_en               ),
  .cpurst_b                     (cpurst_b                    ),
  .da_xx_fwd_data               (da_xx_fwd_data              ),
  .da_xx_fwd_dst_reg            (da_xx_fwd_dst_reg           ),
  .da_xx_fwd_vld                (da_xx_fwd_vld               ),
  .forever_cpuclk               (forever_cpuclk              ),
  .hpcp_iu_cnt_en               (hpcp_iu_cnt_en              ),
  .idu_alu_ex1_gateclk_sel      (idu_alu_ex1_gateclk_sel     ),
  .idu_bju_ex1_gateclk_sel      (idu_bju_ex1_gateclk_sel     ),
  .idu_div_ex1_gateclk_sel      (idu_div_ex1_gateclk_sel     ),
  .idu_iu_ex1_alu_dp_sel        (idu_iu_ex1_alu_dp_sel       ),
  .idu_iu_ex1_alu_sel           (idu_iu_ex1_alu_sel          ),
  .idu_iu_ex1_bht_pred          (idu_iu_ex1_bht_pred         ),
  .idu_iu_ex1_bju_br_sel        (idu_iu_ex1_bju_br_sel       ),
  .idu_iu_ex1_bju_dp_sel        (idu_iu_ex1_bju_dp_sel       ),
  .idu_iu_ex1_bju_sel           (idu_iu_ex1_bju_sel          ),
  .idu_iu_ex1_div_dp_sel        (idu_iu_ex1_div_dp_sel       ),
  .idu_iu_ex1_div_sel           (idu_iu_ex1_div_sel          ),
  .idu_iu_ex1_dst0_reg          (idu_iu_ex1_dst0_reg         ),
  .idu_iu_ex1_func              (idu_iu_ex1_func             ),
  .idu_iu_ex1_inst_vld          (idu_iu_ex1_inst_vld         ),
  .idu_iu_ex1_length            (idu_iu_ex1_length           ),
  .idu_iu_ex1_mult_dp_sel       (idu_iu_ex1_mult_dp_sel      ),
  .idu_iu_ex1_mult_sel          (idu_iu_ex1_mult_sel         ),
  .idu_iu_ex1_pipedown_vld      (idu_iu_ex1_pipedown_vld     ),
  .idu_iu_ex1_split             (idu_iu_ex1_split            ),
  .idu_iu_ex1_src0_data         (idu_iu_ex1_src0_data        ),
  .idu_iu_ex1_src0_ready        (idu_iu_ex1_src0_ready       ),
  .idu_iu_ex1_src0_reg          (idu_iu_ex1_src0_reg         ),
  .idu_iu_ex1_src1_data         (idu_iu_ex1_src1_data        ),
  .idu_iu_ex1_src1_ready        (idu_iu_ex1_src1_ready       ),
  .idu_iu_ex1_src1_reg          (idu_iu_ex1_src1_reg         ),
  .idu_iu_ex1_src2_data         (idu_iu_ex1_src2_data        ),
  .idu_mult_ex1_gateclk_sel     (idu_mult_ex1_gateclk_sel    ),
  .ifu_iu_chgflw_pc             (ifu_iu_chgflw_pc            ),
  .ifu_iu_chgflw_vld            (ifu_iu_chgflw_vld           ),
  .ifu_iu_ex1_pc_pred           (ifu_iu_ex1_pc_pred          ),
  .ifu_iu_reset_vld             (ifu_iu_reset_vld            ),
  .ifu_iu_warm_up               (ifu_iu_warm_up              ),
  .iu_cp0_ex1_cur_pc            (iu_cp0_ex1_cur_pc           ),
  .iu_dtu_debug_info            (iu_dtu_debug_info           ),
  .iu_hpcp_inst_bht_mispred     (iu_hpcp_inst_bht_mispred    ),
  .iu_hpcp_inst_condbr          (iu_hpcp_inst_condbr         ),
  .iu_hpcp_jump_8m              (iu_hpcp_jump_8m             ),
  .iu_idu_bju_full              (iu_idu_bju_full             ),
  .iu_idu_bju_global_full       (iu_idu_bju_global_full      ),
  .iu_idu_div_full              (iu_idu_div_full             ),
  .iu_idu_mult_full             (iu_idu_mult_full            ),
  .iu_idu_mult_issue_stall      (iu_idu_mult_issue_stall     ),
  .iu_ifu_bht_cur_pc            (iu_ifu_bht_cur_pc           ),
  .iu_ifu_bht_mispred           (iu_ifu_bht_mispred          ),
  .iu_ifu_bht_mispred_gate      (iu_ifu_bht_mispred_gate     ),
  .iu_ifu_bht_pred              (iu_ifu_bht_pred             ),
  .iu_ifu_bht_taken             (iu_ifu_bht_taken            ),
  .iu_ifu_br_vld                (iu_ifu_br_vld               ),
  .iu_ifu_br_vld_gate           (iu_ifu_br_vld_gate          ),
  .iu_ifu_link_vld              (iu_ifu_link_vld             ),
  .iu_ifu_link_vld_gate         (iu_ifu_link_vld_gate        ),
  .iu_ifu_pc_mispred            (iu_ifu_pc_mispred           ),
  .iu_ifu_pc_mispred_gate       (iu_ifu_pc_mispred_gate      ),
  .iu_ifu_ret_vld               (iu_ifu_ret_vld              ),
  .iu_ifu_ret_vld_gate          (iu_ifu_ret_vld_gate         ),
  .iu_ifu_tar_pc                (iu_ifu_tar_pc               ),
  .iu_ifu_tar_pc_vld            (iu_ifu_tar_pc_vld           ),
  .iu_ifu_tar_pc_vld_gate       (iu_ifu_tar_pc_vld_gate      ),
  .iu_lsu_ex1_cur_pc            (iu_lsu_ex1_cur_pc           ),
  .iu_rtu_depd_lsu_chgflow_vld  (iu_rtu_depd_lsu_chgflow_vld ),
  .iu_rtu_depd_lsu_next_pc      (iu_rtu_depd_lsu_next_pc     ),
  .iu_rtu_div_data              (iu_rtu_div_data             ),
  .iu_rtu_div_preg              (iu_rtu_div_preg             ),
  .iu_rtu_div_wb_dp             (iu_rtu_div_wb_dp            ),
  .iu_rtu_div_wb_vld            (iu_rtu_div_wb_vld           ),
  .iu_rtu_ex1_alu_cmplt         (iu_rtu_ex1_alu_cmplt        ),
  .iu_rtu_ex1_alu_cmplt_dp      (iu_rtu_ex1_alu_cmplt_dp     ),
  .iu_rtu_ex1_alu_data          (iu_rtu_ex1_alu_data         ),
  .iu_rtu_ex1_alu_inst_len      (iu_rtu_ex1_alu_inst_len     ),
  .iu_rtu_ex1_alu_inst_split    (iu_rtu_ex1_alu_inst_split   ),
  .iu_rtu_ex1_alu_preg          (iu_rtu_ex1_alu_preg         ),
  .iu_rtu_ex1_alu_wb_dp         (iu_rtu_ex1_alu_wb_dp        ),
  .iu_rtu_ex1_alu_wb_vld        (iu_rtu_ex1_alu_wb_vld       ),
  .iu_rtu_ex1_bju_cmplt         (iu_rtu_ex1_bju_cmplt        ),
  .iu_rtu_ex1_bju_cmplt_dp      (iu_rtu_ex1_bju_cmplt_dp     ),
  .iu_rtu_ex1_bju_data          (iu_rtu_ex1_bju_data         ),
  .iu_rtu_ex1_bju_inst_len      (iu_rtu_ex1_bju_inst_len     ),
  .iu_rtu_ex1_bju_preg          (iu_rtu_ex1_bju_preg         ),
  .iu_rtu_ex1_bju_wb_dp         (iu_rtu_ex1_bju_wb_dp        ),
  .iu_rtu_ex1_bju_wb_vld        (iu_rtu_ex1_bju_wb_vld       ),
  .iu_rtu_ex1_branch_inst       (iu_rtu_ex1_branch_inst      ),
  .iu_rtu_ex1_cur_pc            (iu_rtu_ex1_cur_pc           ),
  .iu_rtu_ex1_div_cmplt         (iu_rtu_ex1_div_cmplt        ),
  .iu_rtu_ex1_div_cmplt_dp      (iu_rtu_ex1_div_cmplt_dp     ),
  .iu_rtu_ex1_mul_cmplt         (iu_rtu_ex1_mul_cmplt        ),
  .iu_rtu_ex1_mul_cmplt_dp      (iu_rtu_ex1_mul_cmplt_dp     ),
  .iu_rtu_ex1_next_pc           (iu_rtu_ex1_next_pc          ),
  .iu_rtu_ex2_bju_ras_mispred   (iu_rtu_ex2_bju_ras_mispred  ),
  .iu_rtu_ex3_mul_data          (iu_rtu_ex3_mul_data         ),
  .iu_rtu_ex3_mul_preg          (iu_rtu_ex3_mul_preg         ),
  .iu_rtu_ex3_mul_wb_vld        (iu_rtu_ex3_mul_wb_vld       ),
  .iu_xx_no_op                  (iu_xx_no_op                 ),
  .iu_yy_xx_cancel              (iu_yy_xx_cancel             ),
  .lsu_iu_ex2_data              (lsu_iu_ex2_data             ),
  .lsu_iu_ex2_data_vld          (lsu_iu_ex2_data_vld         ),
  .lsu_iu_ex2_dest_reg          (lsu_iu_ex2_dest_reg         ),
  .mmu_xx_mmu_en                (mmu_xx_mmu_en               ),
  .pad_yy_icg_scan_en           (pad_yy_icg_scan_en          ),
  .rtu_iu_div_wb_grant          (rtu_iu_div_wb_grant         ),
  .rtu_iu_div_wb_grant_for_full (rtu_iu_div_wb_grant_for_full),
  .rtu_iu_ex1_cmplt             (rtu_iu_ex1_cmplt            ),
  .rtu_iu_ex1_cmplt_dp          (rtu_iu_ex1_cmplt_dp         ),
  .rtu_iu_ex1_inst_len          (rtu_iu_ex1_inst_len         ),
  .rtu_iu_ex1_inst_split        (rtu_iu_ex1_inst_split       ),
  .rtu_iu_ex2_cur_pc            (rtu_iu_ex2_cur_pc           ),
  .rtu_iu_ex2_next_pc           (rtu_iu_ex2_next_pc          ),
  .rtu_iu_mul_wb_grant          (rtu_iu_mul_wb_grant         ),
  .rtu_iu_mul_wb_grant_for_full (rtu_iu_mul_wb_grant_for_full),
  .rtu_yy_xx_flush_fe           (rtu_yy_xx_flush_fe          )
);

aq_vpu_top  x_aq_vpu_top (
  .cp0_vpu_icg_en                   (cp0_vpu_icg_en                  ),
  .cp0_vpu_xx_bf16                  (cp0_vpu_xx_bf16                 ),
  .cp0_vpu_xx_dqnan                 (cp0_vpu_xx_dqnan                ),
  .cp0_vpu_xx_rm                    (cp0_vpu_xx_rm                   ),
  .cp0_yy_clk_en                    (cp0_yy_clk_en                   ),
  .cpurst_b                         (cpurst_b                        ),
  .forever_cpuclk                   (forever_cpuclk                  ),
  .ifu_vpu_warm_up                  (ifu_vpu_warm_up                 ),
  .lsu_vlsu_bytes_vld               (lsu_vlsu_bytes_vld              ),
  .lsu_vlsu_data                    (lsu_vlsu_data                   ),
  .lsu_vlsu_data_grant              (lsu_vlsu_data_grant             ),
  .lsu_vlsu_data_vld                (lsu_vlsu_data_vld               ),
  .lsu_vlsu_dc_create_vld           (lsu_vlsu_dc_create_vld          ),
  .lsu_vlsu_dc_fld_req              (lsu_vlsu_dc_fld_req             ),
  .lsu_vlsu_dc_fof                  (lsu_vlsu_dc_fof                 ),
  .lsu_vlsu_dc_nf                   (lsu_vlsu_dc_nf                  ),
  .lsu_vlsu_dc_sew                  (lsu_vlsu_dc_sew                 ),
  .lsu_vlsu_dc_split_cnt            (lsu_vlsu_dc_split_cnt           ),
  .lsu_vlsu_dc_sseg_first           (lsu_vlsu_dc_sseg_first          ),
  .lsu_vlsu_dc_stall                (lsu_vlsu_dc_stall               ),
  .lsu_vlsu_dest_reg                (lsu_vlsu_dest_reg               ),
  .lsu_vlsu_expt_vld                (lsu_vlsu_expt_vld               ),
  .lsu_vlsu_func                    (lsu_vlsu_func                   ),
  .lsu_vlsu_sew                     (lsu_vlsu_sew                    ),
  .lsu_vlsu_split_last              (lsu_vlsu_split_last             ),
  .lsu_vlsu_st_expt                 (lsu_vlsu_st_expt                ),
  .lsu_vlsu_st_offset               (lsu_vlsu_st_offset              ),
  .lsu_vlsu_st_sew                  (lsu_vlsu_st_sew                 ),
  .lsu_vlsu_st_size                 (lsu_vlsu_st_size                ),
  .lsu_vlsu_vl_update               (lsu_vlsu_vl_update              ),
  .lsu_vlsu_vl_upval                (lsu_vlsu_vl_upval               ),
  .pad_yy_icg_scan_en               (pad_yy_icg_scan_en              ),
  .rtu_vpu_gpr_wb_grnt              (rtu_vpu_gpr_wb_grnt             ),
  .rtu_yy_xx_async_flush            (rtu_yy_xx_async_flush           ),
  .rtu_yy_xx_flush                  (rtu_yy_xx_flush                 ),
  .vidu_vpu_vid_fp_inst_dp_vld      (vidu_vpu_vid_fp_inst_dp_vld     ),
  .vidu_vpu_vid_fp_inst_dst_reg     (vidu_vpu_vid_fp_inst_dst_reg    ),
  .vidu_vpu_vid_fp_inst_dst_vld     (vidu_vpu_vid_fp_inst_dst_vld    ),
  .vidu_vpu_vid_fp_inst_dste_vld    (vidu_vpu_vid_fp_inst_dste_vld   ),
  .vidu_vpu_vid_fp_inst_dstf_reg    (vidu_vpu_vid_fp_inst_dstf_reg   ),
  .vidu_vpu_vid_fp_inst_dstf_vld    (vidu_vpu_vid_fp_inst_dstf_vld   ),
  .vidu_vpu_vid_fp_inst_eu          (vidu_vpu_vid_fp_inst_eu         ),
  .vidu_vpu_vid_fp_inst_func        (vidu_vpu_vid_fp_inst_func       ),
  .vidu_vpu_vid_fp_inst_gateclk_vld (vidu_vpu_vid_fp_inst_gateclk_vld),
  .vidu_vpu_vid_fp_inst_src1_data   (vidu_vpu_vid_fp_inst_src1_data  ),
  .vidu_vpu_vid_fp_inst_srcf0_data  (vidu_vpu_vid_fp_inst_srcf0_data ),
  .vidu_vpu_vid_fp_inst_srcf1_data  (vidu_vpu_vid_fp_inst_srcf1_data ),
  .vidu_vpu_vid_fp_inst_srcf2_data  (vidu_vpu_vid_fp_inst_srcf2_data ),
  .vidu_vpu_vid_fp_inst_srcf2_rdy   (vidu_vpu_vid_fp_inst_srcf2_rdy  ),
  .vidu_vpu_vid_fp_inst_srcf2_vld   (vidu_vpu_vid_fp_inst_srcf2_vld  ),
  .vidu_vpu_vid_fp_inst_vld         (vidu_vpu_vid_fp_inst_vld        ),
  .vlsu_buf_stall                   (vlsu_buf_stall                  ),
  .vlsu_dtu_data                    (vlsu_dtu_data                   ),
  .vlsu_dtu_data_vld                (vlsu_dtu_data_vld               ),
  .vlsu_dtu_data_vld_gate           (vlsu_dtu_data_vld_gate          ),
  .vlsu_lsu_data_shift              (vlsu_lsu_data_shift             ),
  .vlsu_lsu_data_vld                (vlsu_lsu_data_vld               ),
  .vlsu_lsu_fwd_data                (vlsu_lsu_fwd_data               ),
  .vlsu_lsu_fwd_dest_reg            (vlsu_lsu_fwd_dest_reg           ),
  .vlsu_lsu_fwd_vld                 (vlsu_lsu_fwd_vld                ),
  .vlsu_lsu_src2_depd               (vlsu_lsu_src2_depd              ),
  .vlsu_lsu_src2_reg                (vlsu_lsu_src2_reg               ),
  .vlsu_lsu_wdata                   (vlsu_lsu_wdata                  ),
  .vlsu_rtu_vl_updt_data            (vlsu_rtu_vl_updt_data           ),
  .vlsu_rtu_vl_updt_vld             (vlsu_rtu_vl_updt_vld            ),
  .vlsu_xx_no_op                    (vlsu_xx_no_op                   ),
  .vpu_dtu_dbg_info                 (vpu_dtu_dbg_info                ),
  .vpu_rtu_fflag                    (vpu_rtu_fflag                   ),
  .vpu_rtu_fflag_vld                (vpu_rtu_fflag_vld               ),
  .vpu_rtu_gpr_wb_data              (vpu_rtu_gpr_wb_data             ),
  .vpu_rtu_gpr_wb_index             (vpu_rtu_gpr_wb_index            ),
  .vpu_rtu_gpr_wb_req               (vpu_rtu_gpr_wb_req              ),
  .vpu_rtu_no_op                    (vpu_rtu_no_op                   ),
  .vpu_vidu_fp_fwd_data             (vpu_vidu_fp_fwd_data            ),
  .vpu_vidu_fp_fwd_reg              (vpu_vidu_fp_fwd_reg             ),
  .vpu_vidu_fp_fwd_vld              (vpu_vidu_fp_fwd_vld             ),
  .vpu_vidu_fp_wb_data              (vpu_vidu_fp_wb_data             ),
  .vpu_vidu_fp_wb_reg               (vpu_vidu_fp_wb_reg              ),
  .vpu_vidu_fp_wb_vld               (vpu_vidu_fp_wb_vld              ),
  .vpu_vidu_vex1_fp_stall           (vpu_vidu_vex1_fp_stall          ),
  .vpu_vidu_wbt_fp_wb0_reg          (vpu_vidu_wbt_fp_wb0_reg         ),
  .vpu_vidu_wbt_fp_wb0_vld          (vpu_vidu_wbt_fp_wb0_vld         ),
  .vpu_vidu_wbt_fp_wb1_reg          (vpu_vidu_wbt_fp_wb1_reg         ),
  .vpu_vidu_wbt_fp_wb1_vld          (vpu_vidu_wbt_fp_wb1_vld         )
);

aq_lsu_top  x_aq_lsu_top (
  .biu_lsu_arready              (biu_lsu_arready             ),
  .biu_lsu_no_op                (biu_lsu_no_op               ),
  .biu_lsu_rdata                (biu_lsu_rdata               ),
  .biu_lsu_rid                  (biu_lsu_rid                 ),
  .biu_lsu_rlast                (biu_lsu_rlast               ),
  .biu_lsu_rresp                (biu_lsu_rresp               ),
  .biu_lsu_rvalid               (biu_lsu_rvalid              ),
  .biu_lsu_stb_awready          (biu_lsu_stb_awready         ),
  .biu_lsu_stb_wready           (biu_lsu_stb_wready          ),
  .biu_lsu_vb_awready           (biu_lsu_vb_awready          ),
  .biu_lsu_vb_wready            (biu_lsu_vb_wready           ),
  .cp0_lsu_amr                  (cp0_lsu_amr                 ),
  .cp0_lsu_dcache_en            (cp0_lsu_dcache_en           ),
  .cp0_lsu_dcache_pref_dist     (cp0_lsu_dcache_pref_dist    ),
  .cp0_lsu_dcache_pref_en       (cp0_lsu_dcache_pref_en      ),
  .cp0_lsu_dcache_read_idx      (cp0_lsu_dcache_read_idx     ),
  .cp0_lsu_dcache_read_req      (cp0_lsu_dcache_read_req     ),
  .cp0_lsu_dcache_read_type     (cp0_lsu_dcache_read_type    ),
  .cp0_lsu_dcache_read_way      (cp0_lsu_dcache_read_way     ),
  .cp0_lsu_dcache_wa            (cp0_lsu_dcache_wa           ),
  .cp0_lsu_dcache_wb            (cp0_lsu_dcache_wb           ),
  .cp0_lsu_fence_req            (cp0_lsu_fence_req           ),
  .cp0_lsu_icc_addr             (cp0_lsu_icc_addr            ),
  .cp0_lsu_icc_op               (cp0_lsu_icc_op              ),
  .cp0_lsu_icc_req              (cp0_lsu_icc_req             ),
  .cp0_lsu_icc_type             (cp0_lsu_icc_type            ),
  .cp0_lsu_icg_en               (cp0_lsu_icg_en              ),
  .cp0_lsu_mm                   (cp0_lsu_mm                  ),
  .cp0_lsu_mpp                  (cp0_lsu_mpp                 ),
  .cp0_lsu_mprv                 (cp0_lsu_mprv                ),
  .cp0_lsu_sync_req             (cp0_lsu_sync_req            ),
  .cp0_lsu_we_en                (cp0_lsu_we_en               ),
  .cp0_yy_priv_mode             (cp0_yy_priv_mode            ),
  .cpurst_b                     (cpurst_b                    ),
  .da_xx_fwd_data               (da_xx_fwd_data              ),
  .da_xx_fwd_dst_reg            (da_xx_fwd_dst_reg           ),
  .da_xx_fwd_vld                (da_xx_fwd_vld               ),
  .dtu_lsu_addr_trig_en         (dtu_lsu_addr_trig_en        ),
  .dtu_lsu_data_trig_en         (dtu_lsu_data_trig_en        ),
  .dtu_lsu_halt_info            (dtu_lsu_halt_info           ),
  .dtu_lsu_halt_info_vld        (dtu_lsu_halt_info_vld       ),
  .forever_cpuclk               (forever_cpuclk              ),
  .hpcp_lsu_cnt_en              (hpcp_lsu_cnt_en             ),
  .idu_lsu_ex1_dp_sel           (idu_lsu_ex1_dp_sel          ),
  .idu_lsu_ex1_dst0_reg         (idu_lsu_ex1_dst0_reg        ),
  .idu_lsu_ex1_dst1_reg         (idu_lsu_ex1_dst1_reg        ),
  .idu_lsu_ex1_func             (idu_lsu_ex1_func            ),
  .idu_lsu_ex1_gateclk_sel      (idu_lsu_ex1_gateclk_sel     ),
  .idu_lsu_ex1_halt_info        (idu_lsu_ex1_halt_info       ),
  .idu_lsu_ex1_length           (idu_lsu_ex1_length          ),
  .idu_lsu_ex1_sel              (idu_lsu_ex1_sel             ),
  .idu_lsu_ex1_split            (idu_lsu_ex1_split           ),
  .idu_lsu_ex1_src0_data        (idu_lsu_ex1_src0_data       ),
  .idu_lsu_ex1_src1_data        (idu_lsu_ex1_src1_data       ),
  .idu_lsu_ex1_src2_data        (idu_lsu_ex1_src2_data       ),
  .idu_lsu_ex1_src2_ready       (idu_lsu_ex1_src2_ready      ),
  .idu_lsu_ex1_src2_reg         (idu_lsu_ex1_src2_reg        ),
  .idu_lsu_ex1_vlmul            (idu_lsu_ex1_vlmul           ),
  .idu_lsu_ex1_vsew             (idu_lsu_ex1_vsew            ),
  .ifu_lsu_warm_up              (ifu_lsu_warm_up             ),
  .iu_lsu_ex1_cur_pc            (iu_lsu_ex1_cur_pc           ),
  .lsu_biu_araddr               (lsu_biu_araddr              ),
  .lsu_biu_arburst              (lsu_biu_arburst             ),
  .lsu_biu_arcache              (lsu_biu_arcache             ),
  .lsu_biu_arid                 (lsu_biu_arid                ),
  .lsu_biu_arlen                (lsu_biu_arlen               ),
  .lsu_biu_arprot               (lsu_biu_arprot              ),
  .lsu_biu_arsize               (lsu_biu_arsize              ),
  .lsu_biu_aruser               (lsu_biu_aruser              ),
  .lsu_biu_arvalid              (lsu_biu_arvalid             ),
  .lsu_biu_stb_awaddr           (lsu_biu_stb_awaddr          ),
  .lsu_biu_stb_awburst          (lsu_biu_stb_awburst         ),
  .lsu_biu_stb_awcache          (lsu_biu_stb_awcache         ),
  .lsu_biu_stb_awid             (lsu_biu_stb_awid            ),
  .lsu_biu_stb_awlen            (lsu_biu_stb_awlen           ),
  .lsu_biu_stb_awprot           (lsu_biu_stb_awprot          ),
  .lsu_biu_stb_awsize           (lsu_biu_stb_awsize          ),
  .lsu_biu_stb_awuser           (lsu_biu_stb_awuser          ),
  .lsu_biu_stb_awvalid          (lsu_biu_stb_awvalid         ),
  .lsu_biu_stb_wdata            (lsu_biu_stb_wdata           ),
  .lsu_biu_stb_wlast            (lsu_biu_stb_wlast           ),
  .lsu_biu_stb_wstrb            (lsu_biu_stb_wstrb           ),
  .lsu_biu_stb_wvalid           (lsu_biu_stb_wvalid          ),
  .lsu_biu_vb_awaddr            (lsu_biu_vb_awaddr           ),
  .lsu_biu_vb_awburst           (lsu_biu_vb_awburst          ),
  .lsu_biu_vb_awcache           (lsu_biu_vb_awcache          ),
  .lsu_biu_vb_awid              (lsu_biu_vb_awid             ),
  .lsu_biu_vb_awlen             (lsu_biu_vb_awlen            ),
  .lsu_biu_vb_awprot            (lsu_biu_vb_awprot           ),
  .lsu_biu_vb_awsize            (lsu_biu_vb_awsize           ),
  .lsu_biu_vb_awvalid           (lsu_biu_vb_awvalid          ),
  .lsu_biu_vb_wdata             (lsu_biu_vb_wdata            ),
  .lsu_biu_vb_wlast             (lsu_biu_vb_wlast            ),
  .lsu_biu_vb_wstrb             (lsu_biu_vb_wstrb            ),
  .lsu_biu_vb_wvalid            (lsu_biu_vb_wvalid           ),
  .lsu_cp0_dcache_read_data     (lsu_cp0_dcache_read_data    ),
  .lsu_cp0_dcache_read_data_vld (lsu_cp0_dcache_read_data_vld),
  .lsu_cp0_fence_ack            (lsu_cp0_fence_ack           ),
  .lsu_cp0_icc_done             (lsu_cp0_icc_done            ),
  .lsu_cp0_sync_ack             (lsu_cp0_sync_ack            ),
  .lsu_dtu_debug_info           (lsu_dtu_debug_info          ),
  .lsu_dtu_halt_info            (lsu_dtu_halt_info           ),
  .lsu_dtu_last_check           (lsu_dtu_last_check          ),
  .lsu_dtu_ldst_addr            (lsu_dtu_ldst_addr           ),
  .lsu_dtu_ldst_addr_vld        (lsu_dtu_ldst_addr_vld       ),
  .lsu_dtu_ldst_bytes_vld       (lsu_dtu_ldst_bytes_vld      ),
  .lsu_dtu_ldst_data            (lsu_dtu_ldst_data           ),
  .lsu_dtu_ldst_data_vld        (lsu_dtu_ldst_data_vld       ),
  .lsu_dtu_ldst_type            (lsu_dtu_ldst_type           ),
  .lsu_dtu_mem_access_size      (lsu_dtu_mem_access_size     ),
  .lsu_hpcp_cache_read_access   (lsu_hpcp_cache_read_access  ),
  .lsu_hpcp_cache_read_miss     (lsu_hpcp_cache_read_miss    ),
  .lsu_hpcp_cache_write_access  (lsu_hpcp_cache_write_access ),
  .lsu_hpcp_cache_write_miss    (lsu_hpcp_cache_write_miss   ),
  .lsu_hpcp_inst_store          (lsu_hpcp_inst_store         ),
  .lsu_hpcp_unalign_inst        (lsu_hpcp_unalign_inst       ),
  .lsu_idu_full                 (lsu_idu_full                ),
  .lsu_idu_global_full          (lsu_idu_global_full         ),
  .lsu_iu_ex2_data              (lsu_iu_ex2_data             ),
  .lsu_iu_ex2_data_vld          (lsu_iu_ex2_data_vld         ),
  .lsu_iu_ex2_dest_reg          (lsu_iu_ex2_dest_reg         ),
  .lsu_mmu_abort                (lsu_mmu_abort               ),
  .lsu_mmu_bus_error            (lsu_mmu_bus_error           ),
  .lsu_mmu_data                 (lsu_mmu_data                ),
  .lsu_mmu_data_vld             (lsu_mmu_data_vld            ),
  .lsu_mmu_priv_mode            (lsu_mmu_priv_mode           ),
  .lsu_mmu_st_inst              (lsu_mmu_st_inst             ),
  .lsu_mmu_va                   (lsu_mmu_va                  ),
  .lsu_mmu_va_vld               (lsu_mmu_va_vld              ),
  .lsu_rtu_async_expt_vld       (lsu_rtu_async_expt_vld      ),
  .lsu_rtu_async_ld_inst        (lsu_rtu_async_ld_inst       ),
  .lsu_rtu_async_tval           (lsu_rtu_async_tval          ),
  .lsu_rtu_ex1_buffer_vld       (lsu_rtu_ex1_buffer_vld      ),
  .lsu_rtu_ex1_cmplt            (lsu_rtu_ex1_cmplt           ),
  .lsu_rtu_ex1_cmplt_dp         (lsu_rtu_ex1_cmplt_dp        ),
  .lsu_rtu_ex1_cmplt_for_pcgen  (lsu_rtu_ex1_cmplt_for_pcgen ),
  .lsu_rtu_ex1_data             (lsu_rtu_ex1_data            ),
  .lsu_rtu_ex1_dest_reg         (lsu_rtu_ex1_dest_reg        ),
  .lsu_rtu_ex1_expt_tval        (lsu_rtu_ex1_expt_tval       ),
  .lsu_rtu_ex1_expt_vec         (lsu_rtu_ex1_expt_vec        ),
  .lsu_rtu_ex1_expt_vld         (lsu_rtu_ex1_expt_vld        ),
  .lsu_rtu_ex1_fs_dirty         (lsu_rtu_ex1_fs_dirty        ),
  .lsu_rtu_ex1_halt_info        (lsu_rtu_ex1_halt_info       ),
  .lsu_rtu_ex1_inst_len         (lsu_rtu_ex1_inst_len        ),
  .lsu_rtu_ex1_inst_split       (lsu_rtu_ex1_inst_split      ),
  .lsu_rtu_ex1_tval2_vld        (lsu_rtu_ex1_tval2_vld       ),
  .lsu_rtu_ex1_vs_dirty         (lsu_rtu_ex1_vs_dirty        ),
  .lsu_rtu_ex1_vstart           (lsu_rtu_ex1_vstart          ),
  .lsu_rtu_ex1_vstart_vld       (lsu_rtu_ex1_vstart_vld      ),
  .lsu_rtu_ex1_wb_dp            (lsu_rtu_ex1_wb_dp           ),
  .lsu_rtu_ex1_wb_vld           (lsu_rtu_ex1_wb_vld          ),
  .lsu_rtu_ex2_data             (lsu_rtu_ex2_data            ),
  .lsu_rtu_ex2_data_vld         (lsu_rtu_ex2_data_vld        ),
  .lsu_rtu_ex2_dest_reg         (lsu_rtu_ex2_dest_reg        ),
  .lsu_rtu_ex2_tval2            (lsu_rtu_ex2_tval2           ),
  .lsu_rtu_no_op                (lsu_rtu_no_op               ),
  .lsu_rtu_wb_data              (lsu_rtu_wb_data             ),
  .lsu_rtu_wb_dest_reg          (lsu_rtu_wb_dest_reg         ),
  .lsu_rtu_wb_vld               (lsu_rtu_wb_vld              ),
  .lsu_vlsu_bytes_vld           (lsu_vlsu_bytes_vld          ),
  .lsu_vlsu_data                (lsu_vlsu_data               ),
  .lsu_vlsu_data_grant          (lsu_vlsu_data_grant         ),
  .lsu_vlsu_data_vld            (lsu_vlsu_data_vld           ),
  .lsu_vlsu_dc_create_vld       (lsu_vlsu_dc_create_vld      ),
  .lsu_vlsu_dc_fld_req          (lsu_vlsu_dc_fld_req         ),
  .lsu_vlsu_dc_fof              (lsu_vlsu_dc_fof             ),
  .lsu_vlsu_dc_nf               (lsu_vlsu_dc_nf              ),
  .lsu_vlsu_dc_sew              (lsu_vlsu_dc_sew             ),
  .lsu_vlsu_dc_split_cnt        (lsu_vlsu_dc_split_cnt       ),
  .lsu_vlsu_dc_sseg_first       (lsu_vlsu_dc_sseg_first      ),
  .lsu_vlsu_dc_stall            (lsu_vlsu_dc_stall           ),
  .lsu_vlsu_dest_reg            (lsu_vlsu_dest_reg           ),
  .lsu_vlsu_expt_vld            (lsu_vlsu_expt_vld           ),
  .lsu_vlsu_func                (lsu_vlsu_func               ),
  .lsu_vlsu_sew                 (lsu_vlsu_sew                ),
  .lsu_vlsu_split_last          (lsu_vlsu_split_last         ),
  .lsu_vlsu_st_expt             (lsu_vlsu_st_expt            ),
  .lsu_vlsu_st_offset           (lsu_vlsu_st_offset          ),
  .lsu_vlsu_st_sew              (lsu_vlsu_st_sew             ),
  .lsu_vlsu_st_size             (lsu_vlsu_st_size            ),
  .lsu_vlsu_vl_update           (lsu_vlsu_vl_update          ),
  .lsu_vlsu_vl_upval            (lsu_vlsu_vl_upval           ),
  .mmu_lsu_access_fault         (mmu_lsu_access_fault        ),
  .mmu_lsu_buf                  (mmu_lsu_buf                 ),
  .mmu_lsu_ca                   (mmu_lsu_ca                  ),
  .mmu_lsu_data_req             (mmu_lsu_data_req            ),
  .mmu_lsu_data_req_addr        (mmu_lsu_data_req_addr       ),
  .mmu_lsu_data_req_size        (mmu_lsu_data_req_size       ),
  .mmu_lsu_pa                   (mmu_lsu_pa                  ),
  .mmu_lsu_pa_vld               (mmu_lsu_pa_vld              ),
  .mmu_lsu_page_fault           (mmu_lsu_page_fault          ),
  .mmu_lsu_sec                  (mmu_lsu_sec                 ),
  .mmu_lsu_sh                   (mmu_lsu_sh                  ),
  .mmu_lsu_so                   (mmu_lsu_so                  ),
  .pad_yy_icg_scan_en           (pad_yy_icg_scan_en          ),
  .rtu_lsu_async_expt_ack       (rtu_lsu_async_expt_ack      ),
  .rtu_lsu_expt_ack             (rtu_lsu_expt_ack            ),
  .rtu_lsu_expt_exit            (rtu_lsu_expt_exit           ),
  .rtu_yy_xx_async_flush        (rtu_yy_xx_async_flush       ),
  .rtu_yy_xx_dbgon              (rtu_yy_xx_dbgon             ),
  .rtu_yy_xx_flush              (rtu_yy_xx_flush             ),
  .vlsu_buf_stall               (vlsu_buf_stall              ),
  .vlsu_dtu_data                (vlsu_dtu_data               ),
  .vlsu_dtu_data_vld            (vlsu_dtu_data_vld           ),
  .vlsu_dtu_data_vld_gate       (vlsu_dtu_data_vld_gate      ),
  .vlsu_lsu_data_shift          (vlsu_lsu_data_shift         ),
  .vlsu_lsu_data_vld            (vlsu_lsu_data_vld           ),
  .vlsu_lsu_fwd_data            (vlsu_lsu_fwd_data           ),
  .vlsu_lsu_fwd_dest_reg        (vlsu_lsu_fwd_dest_reg       ),
  .vlsu_lsu_fwd_vld             (vlsu_lsu_fwd_vld            ),
  .vlsu_lsu_src2_depd           (vlsu_lsu_src2_depd          ),
  .vlsu_lsu_src2_reg            (vlsu_lsu_src2_reg           ),
  .vlsu_lsu_wdata               (vlsu_lsu_wdata              ),
  .vlsu_xx_no_op                (vlsu_xx_no_op               )
);

aq_cp0_top  x_aq_cp0_top (
  .biu_cp0_coreid               (biu_cp0_coreid              ),
  .biu_cp0_me_int               (biu_cp0_me_int              ),
  .biu_cp0_ms_int               (biu_cp0_ms_int              ),
  .biu_cp0_mt_int               (biu_cp0_mt_int              ),
  .biu_cp0_rvba                 (biu_cp0_rvba                ),
  .biu_cp0_se_int               (biu_cp0_se_int              ),
  .biu_cp0_ss_int               (biu_cp0_ss_int              ),
  .biu_cp0_st_int               (biu_cp0_st_int              ),
  .cp0_biu_icg_en               (cp0_biu_icg_en              ),
  .cp0_biu_lpmd_b               (cp0_biu_lpmd_b              ),
  .cp0_dtu_addr                 (cp0_dtu_addr                ),
  .cp0_dtu_debug_info           (cp0_dtu_debug_info          ),
  .cp0_dtu_icg_en               (cp0_dtu_icg_en              ),
  .cp0_dtu_mexpt_vld            (cp0_dtu_mexpt_vld           ),
  .cp0_dtu_pcfifo_frz           (cp0_dtu_pcfifo_frz          ),
  .cp0_dtu_rreg                 (cp0_dtu_rreg                ),
  .cp0_dtu_satp                 (cp0_dtu_satp                ),
  .cp0_dtu_wdata                (cp0_dtu_wdata               ),
  .cp0_dtu_wreg                 (cp0_dtu_wreg                ),
  .cp0_hpcp_icg_en              (cp0_hpcp_icg_en             ),
  .cp0_hpcp_index               (cp0_hpcp_index              ),
  .cp0_hpcp_int_off_vld         (cp0_hpcp_int_off_vld        ),
  .cp0_hpcp_mcntwen             (cp0_hpcp_mcntwen            ),
  .cp0_hpcp_pmdm                (cp0_hpcp_pmdm               ),
  .cp0_hpcp_pmds                (cp0_hpcp_pmds               ),
  .cp0_hpcp_pmdu                (cp0_hpcp_pmdu               ),
  .cp0_hpcp_sync_stall_vld      (cp0_hpcp_sync_stall_vld     ),
  .cp0_hpcp_wdata               (cp0_hpcp_wdata              ),
  .cp0_hpcp_wreg                (cp0_hpcp_wreg               ),
  .cp0_idu_cskyee               (cp0_idu_cskyee              ),
  .cp0_idu_dis_fence_in_dbg     (cp0_idu_dis_fence_in_dbg    ),
  .cp0_idu_frm                  (cp0_idu_frm                 ),
  .cp0_idu_fs                   (cp0_idu_fs                  ),
  .cp0_idu_icg_en               (cp0_idu_icg_en              ),
  .cp0_idu_issue_stall          (cp0_idu_issue_stall         ),
  .cp0_idu_ucme                 (cp0_idu_ucme                ),
  .cp0_idu_vill                 (cp0_idu_vill                ),
  .cp0_idu_vl_zero              (cp0_idu_vl_zero             ),
  .cp0_idu_vlmul                (cp0_idu_vlmul               ),
  .cp0_idu_vs                   (cp0_idu_vs                  ),
  .cp0_idu_vsetvl_dis_stall     (cp0_idu_vsetvl_dis_stall    ),
  .cp0_idu_vsew                 (cp0_idu_vsew                ),
  .cp0_idu_vstart               (cp0_idu_vstart              ),
  .cp0_ifu_bht_en               (cp0_ifu_bht_en              ),
  .cp0_ifu_bht_inv              (cp0_ifu_bht_inv             ),
  .cp0_ifu_btb_clr              (cp0_ifu_btb_clr             ),
  .cp0_ifu_btb_en               (cp0_ifu_btb_en              ),
  .cp0_ifu_icache_en            (cp0_ifu_icache_en           ),
  .cp0_ifu_icache_inv_addr      (cp0_ifu_icache_inv_addr     ),
  .cp0_ifu_icache_inv_req       (cp0_ifu_icache_inv_req      ),
  .cp0_ifu_icache_inv_type      (cp0_ifu_icache_inv_type     ),
  .cp0_ifu_icache_pref_en       (cp0_ifu_icache_pref_en      ),
  .cp0_ifu_icache_read_index    (cp0_ifu_icache_read_index   ),
  .cp0_ifu_icache_read_req      (cp0_ifu_icache_read_req     ),
  .cp0_ifu_icache_read_tag      (cp0_ifu_icache_read_tag     ),
  .cp0_ifu_icache_read_way      (cp0_ifu_icache_read_way     ),
  .cp0_ifu_icg_en               (cp0_ifu_icg_en              ),
  .cp0_ifu_in_lpmd              (cp0_ifu_in_lpmd             ),
  .cp0_ifu_iwpe                 (cp0_ifu_iwpe                ),
  .cp0_ifu_lpmd_req             (cp0_ifu_lpmd_req            ),
  .cp0_ifu_ras_en               (cp0_ifu_ras_en              ),
  .cp0_ifu_rst_inv_done         (cp0_ifu_rst_inv_done        ),
  .cp0_iu_icg_en                (cp0_iu_icg_en               ),
  .cp0_lsu_amr                  (cp0_lsu_amr                 ),
  .cp0_lsu_dcache_en            (cp0_lsu_dcache_en           ),
  .cp0_lsu_dcache_pref_dist     (cp0_lsu_dcache_pref_dist    ),
  .cp0_lsu_dcache_pref_en       (cp0_lsu_dcache_pref_en      ),
  .cp0_lsu_dcache_read_idx      (cp0_lsu_dcache_read_idx     ),
  .cp0_lsu_dcache_read_req      (cp0_lsu_dcache_read_req     ),
  .cp0_lsu_dcache_read_type     (cp0_lsu_dcache_read_type    ),
  .cp0_lsu_dcache_read_way      (cp0_lsu_dcache_read_way     ),
  .cp0_lsu_dcache_wa            (cp0_lsu_dcache_wa           ),
  .cp0_lsu_dcache_wb            (cp0_lsu_dcache_wb           ),
  .cp0_lsu_fence_req            (cp0_lsu_fence_req           ),
  .cp0_lsu_icc_addr             (cp0_lsu_icc_addr            ),
  .cp0_lsu_icc_op               (cp0_lsu_icc_op              ),
  .cp0_lsu_icc_req              (cp0_lsu_icc_req             ),
  .cp0_lsu_icc_type             (cp0_lsu_icc_type            ),
  .cp0_lsu_icg_en               (cp0_lsu_icg_en              ),
  .cp0_lsu_mm                   (cp0_lsu_mm                  ),
  .cp0_lsu_mpp                  (cp0_lsu_mpp                 ),
  .cp0_lsu_mprv                 (cp0_lsu_mprv                ),
  .cp0_lsu_sync_req             (cp0_lsu_sync_req            ),
  .cp0_lsu_we_en                (cp0_lsu_we_en               ),
  .cp0_mmu_addr                 (cp0_mmu_addr                ),
  .cp0_mmu_icg_en               (cp0_mmu_icg_en              ),
  .cp0_mmu_lpmd_req             (cp0_mmu_lpmd_req            ),
  .cp0_mmu_maee                 (cp0_mmu_maee                ),
  .cp0_mmu_mxr                  (cp0_mmu_mxr                 ),
  .cp0_mmu_ptw_en               (cp0_mmu_ptw_en              ),
  .cp0_mmu_satp_data            (cp0_mmu_satp_data           ),
  .cp0_mmu_satp_wen             (cp0_mmu_satp_wen            ),
  .cp0_mmu_sum                  (cp0_mmu_sum                 ),
  .cp0_mmu_tlb_all_inv          (cp0_mmu_tlb_all_inv         ),
  .cp0_mmu_tlb_asid             (cp0_mmu_tlb_asid            ),
  .cp0_mmu_tlb_asid_all_inv     (cp0_mmu_tlb_asid_all_inv    ),
  .cp0_mmu_tlb_va               (cp0_mmu_tlb_va              ),
  .cp0_mmu_tlb_va_all_inv       (cp0_mmu_tlb_va_all_inv      ),
  .cp0_mmu_tlb_va_asid_inv      (cp0_mmu_tlb_va_asid_inv     ),
  .cp0_mmu_wdata                (cp0_mmu_wdata               ),
  .cp0_mmu_wreg                 (cp0_mmu_wreg                ),
  .cp0_pmp_addr                 (cp0_pmp_addr                ),
  .cp0_pmp_icg_en               (cp0_pmp_icg_en              ),
  .cp0_pmp_wdata                (cp0_pmp_wdata               ),
  .cp0_pmp_wreg                 (cp0_pmp_wreg                ),
  .cp0_rtu_ex1_chgflw           (cp0_rtu_ex1_chgflw          ),
  .cp0_rtu_ex1_chgflw_pc        (cp0_rtu_ex1_chgflw_pc       ),
  .cp0_rtu_ex1_cmplt            (cp0_rtu_ex1_cmplt           ),
  .cp0_rtu_ex1_cmplt_dp         (cp0_rtu_ex1_cmplt_dp        ),
  .cp0_rtu_ex1_expt_tval        (cp0_rtu_ex1_expt_tval       ),
  .cp0_rtu_ex1_expt_vec         (cp0_rtu_ex1_expt_vec        ),
  .cp0_rtu_ex1_expt_vld         (cp0_rtu_ex1_expt_vld        ),
  .cp0_rtu_ex1_flush            (cp0_rtu_ex1_flush           ),
  .cp0_rtu_ex1_halt_info        (cp0_rtu_ex1_halt_info       ),
  .cp0_rtu_ex1_inst_dret        (cp0_rtu_ex1_inst_dret       ),
  .cp0_rtu_ex1_inst_ebreak      (cp0_rtu_ex1_inst_ebreak     ),
  .cp0_rtu_ex1_inst_len         (cp0_rtu_ex1_inst_len        ),
  .cp0_rtu_ex1_inst_mret        (cp0_rtu_ex1_inst_mret       ),
  .cp0_rtu_ex1_inst_split       (cp0_rtu_ex1_inst_split      ),
  .cp0_rtu_ex1_inst_sret        (cp0_rtu_ex1_inst_sret       ),
  .cp0_rtu_ex1_vs_dirty         (cp0_rtu_ex1_vs_dirty        ),
  .cp0_rtu_ex1_vs_dirty_dp      (cp0_rtu_ex1_vs_dirty_dp     ),
  .cp0_rtu_ex1_wb_data          (cp0_rtu_ex1_wb_data         ),
  .cp0_rtu_ex1_wb_dp            (cp0_rtu_ex1_wb_dp           ),
  .cp0_rtu_ex1_wb_preg          (cp0_rtu_ex1_wb_preg         ),
  .cp0_rtu_ex1_wb_vld           (cp0_rtu_ex1_wb_vld          ),
  .cp0_rtu_fence_idle           (cp0_rtu_fence_idle          ),
  .cp0_rtu_icg_en               (cp0_rtu_icg_en              ),
  .cp0_rtu_in_lpmd              (cp0_rtu_in_lpmd             ),
  .cp0_rtu_int_vld              (cp0_rtu_int_vld             ),
  .cp0_rtu_trap_pc              (cp0_rtu_trap_pc             ),
  .cp0_rtu_vstart_eq_0          (cp0_rtu_vstart_eq_0         ),
  .cp0_vpu_icg_en               (cp0_vpu_icg_en              ),
  .cp0_vpu_xx_bf16              (cp0_vpu_xx_bf16             ),
  .cp0_vpu_xx_dqnan             (cp0_vpu_xx_dqnan            ),
  .cp0_vpu_xx_rm                (cp0_vpu_xx_rm               ),
  .cp0_xx_mrvbr                 (cp0_xx_mrvbr                ),
  .cp0_yy_clk_en                (cp0_yy_clk_en               ),
  .cp0_yy_priv_mode             (cp0_yy_priv_mode            ),
  .cpurst_b                     (cpurst_b                    ),
  .dtu_cp0_dcsr_mprven          (dtu_cp0_dcsr_mprven         ),
  .dtu_cp0_dcsr_prv             (dtu_cp0_dcsr_prv            ),
  .dtu_cp0_rdata                (dtu_cp0_rdata               ),
  .dtu_cp0_wake_up              (dtu_cp0_wake_up             ),
  .forever_cpuclk               (forever_cpuclk              ),
  .hpcp_cp0_data                (hpcp_cp0_data               ),
  .hpcp_cp0_int_vld             (hpcp_cp0_int_vld            ),
  .hpcp_cp0_sce                 (hpcp_cp0_sce                ),
  .idu_cp0_ex1_dp_sel           (idu_cp0_ex1_dp_sel          ),
  .idu_cp0_ex1_dst0_reg         (idu_cp0_ex1_dst0_reg        ),
  .idu_cp0_ex1_expt_acc_error   (idu_cp0_ex1_expt_acc_error  ),
  .idu_cp0_ex1_expt_high        (idu_cp0_ex1_expt_high       ),
  .idu_cp0_ex1_expt_illegal     (idu_cp0_ex1_expt_illegal    ),
  .idu_cp0_ex1_expt_page_fault  (idu_cp0_ex1_expt_page_fault ),
  .idu_cp0_ex1_func             (idu_cp0_ex1_func            ),
  .idu_cp0_ex1_gateclk_sel      (idu_cp0_ex1_gateclk_sel     ),
  .idu_cp0_ex1_halt_info        (idu_cp0_ex1_halt_info       ),
  .idu_cp0_ex1_length           (idu_cp0_ex1_length          ),
  .idu_cp0_ex1_opcode           (idu_cp0_ex1_opcode          ),
  .idu_cp0_ex1_sel              (idu_cp0_ex1_sel             ),
  .idu_cp0_ex1_split            (idu_cp0_ex1_split           ),
  .idu_cp0_ex1_src0_data        (idu_cp0_ex1_src0_data       ),
  .idu_cp0_ex1_src1_data        (idu_cp0_ex1_src1_data       ),
  .ifu_cp0_bht_inv_done         (ifu_cp0_bht_inv_done        ),
  .ifu_cp0_icache_inv_done      (ifu_cp0_icache_inv_done     ),
  .ifu_cp0_icache_read_data     (ifu_cp0_icache_read_data    ),
  .ifu_cp0_icache_read_data_vld (ifu_cp0_icache_read_data_vld),
  .ifu_cp0_rst_inv_req          (ifu_cp0_rst_inv_req         ),
  .ifu_cp0_warm_up              (ifu_cp0_warm_up             ),
  .ifu_yy_xx_no_op              (ifu_yy_xx_no_op             ),
  .iu_cp0_ex1_cur_pc            (iu_cp0_ex1_cur_pc           ),
  .lsu_cp0_dcache_read_data     (lsu_cp0_dcache_read_data    ),
  .lsu_cp0_dcache_read_data_vld (lsu_cp0_dcache_read_data_vld),
  .lsu_cp0_fence_ack            (lsu_cp0_fence_ack           ),
  .lsu_cp0_icc_done             (lsu_cp0_icc_done            ),
  .lsu_cp0_sync_ack             (lsu_cp0_sync_ack            ),
  .mmu_cp0_cmplt                (mmu_cp0_cmplt               ),
  .mmu_cp0_data                 (mmu_cp0_data                ),
  .mmu_cp0_tlb_inv_done         (mmu_cp0_tlb_inv_done        ),
  .mmu_yy_xx_no_op              (mmu_yy_xx_no_op             ),
  .pad_yy_icg_scan_en           (pad_yy_icg_scan_en          ),
  .pmp_cp0_data                 (pmp_cp0_data                ),
  .rtu_cp0_epc                  (rtu_cp0_epc                 ),
  .rtu_cp0_exit_debug           (rtu_cp0_exit_debug          ),
  .rtu_cp0_fflags               (rtu_cp0_fflags              ),
  .rtu_cp0_fflags_updt          (rtu_cp0_fflags_updt         ),
  .rtu_cp0_fs_dirty_updt        (rtu_cp0_fs_dirty_updt       ),
  .rtu_cp0_fs_dirty_updt_dp     (rtu_cp0_fs_dirty_updt_dp    ),
  .rtu_cp0_tval                 (rtu_cp0_tval                ),
  .rtu_cp0_vl                   (rtu_cp0_vl                  ),
  .rtu_cp0_vl_vld               (rtu_cp0_vl_vld              ),
  .rtu_cp0_vs_dirty_updt        (rtu_cp0_vs_dirty_updt       ),
  .rtu_cp0_vs_dirty_updt_dp     (rtu_cp0_vs_dirty_updt_dp    ),
  .rtu_cp0_vstart               (rtu_cp0_vstart              ),
  .rtu_cp0_vstart_vld           (rtu_cp0_vstart_vld          ),
  .rtu_cp0_vxsat                (rtu_cp0_vxsat               ),
  .rtu_cp0_vxsat_vld            (rtu_cp0_vxsat_vld           ),
  .rtu_yy_xx_dbgon              (rtu_yy_xx_dbgon             ),
  .rtu_yy_xx_expt_int           (rtu_yy_xx_expt_int          ),
  .rtu_yy_xx_expt_vec           (rtu_yy_xx_expt_vec          ),
  .rtu_yy_xx_expt_vld           (rtu_yy_xx_expt_vld          ),
  .rtu_yy_xx_flush              (rtu_yy_xx_flush             ),
  .sysio_cp0_apb_base           (sysio_cp0_apb_base          ),
  .vidu_cp0_vid_fof_vld         (vidu_cp0_vid_fof_vld        )
);

aq_rtu_top  x_aq_rtu_top (
  .cp0_rtu_ex1_chgflw            (cp0_rtu_ex1_chgflw           ),
  .cp0_rtu_ex1_chgflw_pc         (cp0_rtu_ex1_chgflw_pc        ),
  .cp0_rtu_ex1_cmplt             (cp0_rtu_ex1_cmplt            ),
  .cp0_rtu_ex1_cmplt_dp          (cp0_rtu_ex1_cmplt_dp         ),
  .cp0_rtu_ex1_expt_tval         (cp0_rtu_ex1_expt_tval        ),
  .cp0_rtu_ex1_expt_vec          (cp0_rtu_ex1_expt_vec         ),
  .cp0_rtu_ex1_expt_vld          (cp0_rtu_ex1_expt_vld         ),
  .cp0_rtu_ex1_flush             (cp0_rtu_ex1_flush            ),
  .cp0_rtu_ex1_halt_info         (cp0_rtu_ex1_halt_info        ),
  .cp0_rtu_ex1_inst_dret         (cp0_rtu_ex1_inst_dret        ),
  .cp0_rtu_ex1_inst_ebreak       (cp0_rtu_ex1_inst_ebreak      ),
  .cp0_rtu_ex1_inst_len          (cp0_rtu_ex1_inst_len         ),
  .cp0_rtu_ex1_inst_mret         (cp0_rtu_ex1_inst_mret        ),
  .cp0_rtu_ex1_inst_split        (cp0_rtu_ex1_inst_split       ),
  .cp0_rtu_ex1_inst_sret         (cp0_rtu_ex1_inst_sret        ),
  .cp0_rtu_ex1_vs_dirty          (cp0_rtu_ex1_vs_dirty         ),
  .cp0_rtu_ex1_vs_dirty_dp       (cp0_rtu_ex1_vs_dirty_dp      ),
  .cp0_rtu_ex1_wb_data           (cp0_rtu_ex1_wb_data          ),
  .cp0_rtu_ex1_wb_dp             (cp0_rtu_ex1_wb_dp            ),
  .cp0_rtu_ex1_wb_preg           (cp0_rtu_ex1_wb_preg          ),
  .cp0_rtu_ex1_wb_vld            (cp0_rtu_ex1_wb_vld           ),
  .cp0_rtu_fence_idle            (cp0_rtu_fence_idle           ),
  .cp0_rtu_icg_en                (cp0_rtu_icg_en               ),
  .cp0_rtu_in_lpmd               (cp0_rtu_in_lpmd              ),
  .cp0_rtu_int_vld               (cp0_rtu_int_vld              ),
  .cp0_rtu_trap_pc               (cp0_rtu_trap_pc              ),
  .cp0_rtu_vstart_eq_0           (cp0_rtu_vstart_eq_0          ),
  .cp0_yy_clk_en                 (cp0_yy_clk_en                ),
  .cpurst_b                      (cpurst_b                     ),
  .dtu_rtu_async_halt_req        (dtu_rtu_async_halt_req       ),
  .dtu_rtu_dpc                   (dtu_rtu_dpc                  ),
  .dtu_rtu_ebreak_action         (dtu_rtu_ebreak_action        ),
  .dtu_rtu_int_mask              (dtu_rtu_int_mask             ),
  .dtu_rtu_pending_tval          (dtu_rtu_pending_tval         ),
  .dtu_rtu_resume_req            (dtu_rtu_resume_req           ),
  .dtu_rtu_step_en               (dtu_rtu_step_en              ),
  .dtu_rtu_sync_flush            (dtu_rtu_sync_flush           ),
  .dtu_rtu_sync_halt_req         (dtu_rtu_sync_halt_req        ),
  .forever_cpuclk                (forever_cpuclk               ),
  .hpcp_rtu_cnt_en               (hpcp_rtu_cnt_en              ),
  .ifu_rtu_reset_halt_req        (ifu_rtu_reset_halt_req       ),
  .ifu_rtu_warm_up               (ifu_rtu_warm_up              ),
  .iu_rtu_depd_lsu_chgflow_vld   (iu_rtu_depd_lsu_chgflow_vld  ),
  .iu_rtu_depd_lsu_next_pc       (iu_rtu_depd_lsu_next_pc      ),
  .iu_rtu_div_data               (iu_rtu_div_data              ),
  .iu_rtu_div_preg               (iu_rtu_div_preg              ),
  .iu_rtu_div_wb_dp              (iu_rtu_div_wb_dp             ),
  .iu_rtu_div_wb_vld             (iu_rtu_div_wb_vld            ),
  .iu_rtu_ex1_alu_cmplt          (iu_rtu_ex1_alu_cmplt         ),
  .iu_rtu_ex1_alu_cmplt_dp       (iu_rtu_ex1_alu_cmplt_dp      ),
  .iu_rtu_ex1_alu_data           (iu_rtu_ex1_alu_data          ),
  .iu_rtu_ex1_alu_inst_len       (iu_rtu_ex1_alu_inst_len      ),
  .iu_rtu_ex1_alu_inst_split     (iu_rtu_ex1_alu_inst_split    ),
  .iu_rtu_ex1_alu_preg           (iu_rtu_ex1_alu_preg          ),
  .iu_rtu_ex1_alu_wb_dp          (iu_rtu_ex1_alu_wb_dp         ),
  .iu_rtu_ex1_alu_wb_vld         (iu_rtu_ex1_alu_wb_vld        ),
  .iu_rtu_ex1_bju_cmplt          (iu_rtu_ex1_bju_cmplt         ),
  .iu_rtu_ex1_bju_cmplt_dp       (iu_rtu_ex1_bju_cmplt_dp      ),
  .iu_rtu_ex1_bju_data           (iu_rtu_ex1_bju_data          ),
  .iu_rtu_ex1_bju_inst_len       (iu_rtu_ex1_bju_inst_len      ),
  .iu_rtu_ex1_bju_preg           (iu_rtu_ex1_bju_preg          ),
  .iu_rtu_ex1_bju_wb_dp          (iu_rtu_ex1_bju_wb_dp         ),
  .iu_rtu_ex1_bju_wb_vld         (iu_rtu_ex1_bju_wb_vld        ),
  .iu_rtu_ex1_branch_inst        (iu_rtu_ex1_branch_inst       ),
  .iu_rtu_ex1_cur_pc             (iu_rtu_ex1_cur_pc            ),
  .iu_rtu_ex1_div_cmplt          (iu_rtu_ex1_div_cmplt         ),
  .iu_rtu_ex1_div_cmplt_dp       (iu_rtu_ex1_div_cmplt_dp      ),
  .iu_rtu_ex1_mul_cmplt          (iu_rtu_ex1_mul_cmplt         ),
  .iu_rtu_ex1_mul_cmplt_dp       (iu_rtu_ex1_mul_cmplt_dp      ),
  .iu_rtu_ex1_next_pc            (iu_rtu_ex1_next_pc           ),
  .iu_rtu_ex2_bju_ras_mispred    (iu_rtu_ex2_bju_ras_mispred   ),
  .iu_rtu_ex3_mul_data           (iu_rtu_ex3_mul_data          ),
  .iu_rtu_ex3_mul_preg           (iu_rtu_ex3_mul_preg          ),
  .iu_rtu_ex3_mul_wb_vld         (iu_rtu_ex3_mul_wb_vld        ),
  .iu_xx_no_op                   (iu_xx_no_op                  ),
  .lsu_rtu_async_expt_vld        (lsu_rtu_async_expt_vld       ),
  .lsu_rtu_async_ld_inst         (lsu_rtu_async_ld_inst        ),
  .lsu_rtu_async_tval            (lsu_rtu_async_tval           ),
  .lsu_rtu_ex1_buffer_vld        (lsu_rtu_ex1_buffer_vld       ),
  .lsu_rtu_ex1_cmplt             (lsu_rtu_ex1_cmplt            ),
  .lsu_rtu_ex1_cmplt_dp          (lsu_rtu_ex1_cmplt_dp         ),
  .lsu_rtu_ex1_cmplt_for_pcgen   (lsu_rtu_ex1_cmplt_for_pcgen  ),
  .lsu_rtu_ex1_data              (lsu_rtu_ex1_data             ),
  .lsu_rtu_ex1_dest_reg          (lsu_rtu_ex1_dest_reg         ),
  .lsu_rtu_ex1_expt_tval         (lsu_rtu_ex1_expt_tval        ),
  .lsu_rtu_ex1_expt_vec          (lsu_rtu_ex1_expt_vec         ),
  .lsu_rtu_ex1_expt_vld          (lsu_rtu_ex1_expt_vld         ),
  .lsu_rtu_ex1_fs_dirty          (lsu_rtu_ex1_fs_dirty         ),
  .lsu_rtu_ex1_halt_info         (lsu_rtu_ex1_halt_info        ),
  .lsu_rtu_ex1_inst_len          (lsu_rtu_ex1_inst_len         ),
  .lsu_rtu_ex1_inst_split        (lsu_rtu_ex1_inst_split       ),
  .lsu_rtu_ex1_tval2_vld         (lsu_rtu_ex1_tval2_vld        ),
  .lsu_rtu_ex1_vs_dirty          (lsu_rtu_ex1_vs_dirty         ),
  .lsu_rtu_ex1_vstart            (lsu_rtu_ex1_vstart           ),
  .lsu_rtu_ex1_vstart_vld        (lsu_rtu_ex1_vstart_vld       ),
  .lsu_rtu_ex1_wb_dp             (lsu_rtu_ex1_wb_dp            ),
  .lsu_rtu_ex1_wb_vld            (lsu_rtu_ex1_wb_vld           ),
  .lsu_rtu_ex2_data              (lsu_rtu_ex2_data             ),
  .lsu_rtu_ex2_data_vld          (lsu_rtu_ex2_data_vld         ),
  .lsu_rtu_ex2_dest_reg          (lsu_rtu_ex2_dest_reg         ),
  .lsu_rtu_ex2_tval2             (lsu_rtu_ex2_tval2            ),
  .lsu_rtu_no_op                 (lsu_rtu_no_op                ),
  .lsu_rtu_wb_data               (lsu_rtu_wb_data              ),
  .lsu_rtu_wb_dest_reg           (lsu_rtu_wb_dest_reg          ),
  .lsu_rtu_wb_vld                (lsu_rtu_wb_vld               ),
  .mmu_xx_mmu_en                 (mmu_xx_mmu_en                ),
  .pad_yy_icg_scan_en            (pad_yy_icg_scan_en           ),
  .rtu_cp0_epc                   (rtu_cp0_epc                  ),
  .rtu_cp0_exit_debug            (rtu_cp0_exit_debug           ),
  .rtu_cp0_fflags                (rtu_cp0_fflags               ),
  .rtu_cp0_fflags_updt           (rtu_cp0_fflags_updt          ),
  .rtu_cp0_fs_dirty_updt         (rtu_cp0_fs_dirty_updt        ),
  .rtu_cp0_fs_dirty_updt_dp      (rtu_cp0_fs_dirty_updt_dp     ),
  .rtu_cp0_tval                  (rtu_cp0_tval                 ),
  .rtu_cp0_vl                    (rtu_cp0_vl                   ),
  .rtu_cp0_vl_vld                (rtu_cp0_vl_vld               ),
  .rtu_cp0_vs_dirty_updt         (rtu_cp0_vs_dirty_updt        ),
  .rtu_cp0_vs_dirty_updt_dp      (rtu_cp0_vs_dirty_updt_dp     ),
  .rtu_cp0_vstart                (rtu_cp0_vstart               ),
  .rtu_cp0_vstart_vld            (rtu_cp0_vstart_vld           ),
  .rtu_cp0_vxsat                 (rtu_cp0_vxsat                ),
  .rtu_cp0_vxsat_vld             (rtu_cp0_vxsat_vld            ),
  .rtu_cpu_no_retire             (rtu_cpu_no_retire            ),
  .rtu_dtu_debug_info            (rtu_dtu_debug_info           ),
  .rtu_dtu_dpc                   (rtu_dtu_dpc                  ),
  .rtu_dtu_halt_ack              (rtu_dtu_halt_ack             ),
  .rtu_dtu_pending_ack           (rtu_dtu_pending_ack          ),
  .rtu_dtu_retire_chgflw         (rtu_dtu_retire_chgflw        ),
  .rtu_dtu_retire_debug_expt_vld (rtu_dtu_retire_debug_expt_vld),
  .rtu_dtu_retire_halt_info      (rtu_dtu_retire_halt_info     ),
  .rtu_dtu_retire_mret           (rtu_dtu_retire_mret          ),
  .rtu_dtu_retire_next_pc        (rtu_dtu_retire_next_pc       ),
  .rtu_dtu_retire_sret           (rtu_dtu_retire_sret          ),
  .rtu_dtu_retire_vld            (rtu_dtu_retire_vld           ),
  .rtu_dtu_tval                  (rtu_dtu_tval                 ),
  .rtu_hpcp_int_vld              (rtu_hpcp_int_vld             ),
  .rtu_hpcp_retire_inst_vld      (rtu_hpcp_retire_inst_vld     ),
  .rtu_hpcp_retire_pc            (rtu_hpcp_retire_pc           ),
  .rtu_idu_commit                (rtu_idu_commit               ),
  .rtu_idu_commit_for_bju        (rtu_idu_commit_for_bju       ),
  .rtu_idu_flush_fe              (rtu_idu_flush_fe             ),
  .rtu_idu_flush_stall           (rtu_idu_flush_stall          ),
  .rtu_idu_flush_wbt             (rtu_idu_flush_wbt            ),
  .rtu_idu_fwd0_data             (rtu_idu_fwd0_data            ),
  .rtu_idu_fwd0_reg              (rtu_idu_fwd0_reg             ),
  .rtu_idu_fwd0_vld              (rtu_idu_fwd0_vld             ),
  .rtu_idu_fwd1_data             (rtu_idu_fwd1_data            ),
  .rtu_idu_fwd1_reg              (rtu_idu_fwd1_reg             ),
  .rtu_idu_fwd1_vld              (rtu_idu_fwd1_vld             ),
  .rtu_idu_fwd2_data             (rtu_idu_fwd2_data            ),
  .rtu_idu_fwd2_reg              (rtu_idu_fwd2_reg             ),
  .rtu_idu_fwd2_vld              (rtu_idu_fwd2_vld             ),
  .rtu_idu_pipeline_empty        (rtu_idu_pipeline_empty       ),
  .rtu_idu_wb0_data              (rtu_idu_wb0_data             ),
  .rtu_idu_wb0_reg               (rtu_idu_wb0_reg              ),
  .rtu_idu_wb0_vld               (rtu_idu_wb0_vld              ),
  .rtu_idu_wb1_data              (rtu_idu_wb1_data             ),
  .rtu_idu_wb1_reg               (rtu_idu_wb1_reg              ),
  .rtu_idu_wb1_vld               (rtu_idu_wb1_vld              ),
  .rtu_ifu_chgflw_pc             (rtu_ifu_chgflw_pc            ),
  .rtu_ifu_chgflw_vld            (rtu_ifu_chgflw_vld           ),
  .rtu_ifu_dbg_mask              (rtu_ifu_dbg_mask             ),
  .rtu_ifu_flush_fe              (rtu_ifu_flush_fe             ),
  .rtu_iu_div_wb_grant           (rtu_iu_div_wb_grant          ),
  .rtu_iu_div_wb_grant_for_full  (rtu_iu_div_wb_grant_for_full ),
  .rtu_iu_ex1_cmplt              (rtu_iu_ex1_cmplt             ),
  .rtu_iu_ex1_cmplt_dp           (rtu_iu_ex1_cmplt_dp          ),
  .rtu_iu_ex1_inst_len           (rtu_iu_ex1_inst_len          ),
  .rtu_iu_ex1_inst_split         (rtu_iu_ex1_inst_split        ),
  .rtu_iu_ex2_cur_pc             (rtu_iu_ex2_cur_pc            ),
  .rtu_iu_ex2_next_pc            (rtu_iu_ex2_next_pc           ),
  .rtu_iu_mul_wb_grant           (rtu_iu_mul_wb_grant          ),
  .rtu_iu_mul_wb_grant_for_full  (rtu_iu_mul_wb_grant_for_full ),
  .rtu_lsu_async_expt_ack        (rtu_lsu_async_expt_ack       ),
  .rtu_lsu_expt_ack              (rtu_lsu_expt_ack             ),
  .rtu_lsu_expt_exit             (rtu_lsu_expt_exit            ),
  .rtu_mmu_bad_vpn               (rtu_mmu_bad_vpn              ),
  .rtu_mmu_expt_vld              (rtu_mmu_expt_vld             ),
  .rtu_pad_halted                (rtu_pad_halted               ),
  .rtu_pad_retire                (rtu_pad_retire               ),
  .rtu_pad_retire_pc             (rtu_pad_retire_pc            ),
  .rtu_vidu_flush_wbt            (rtu_vidu_flush_wbt           ),
  .rtu_vpu_gpr_wb_grnt           (rtu_vpu_gpr_wb_grnt          ),
  .rtu_yy_xx_async_flush         (rtu_yy_xx_async_flush        ),
  .rtu_yy_xx_dbgon               (rtu_yy_xx_dbgon              ),
  .rtu_yy_xx_expt_int            (rtu_yy_xx_expt_int           ),
  .rtu_yy_xx_expt_vec            (rtu_yy_xx_expt_vec           ),
  .rtu_yy_xx_expt_vld            (rtu_yy_xx_expt_vld           ),
  .rtu_yy_xx_flush               (rtu_yy_xx_flush              ),
  .rtu_yy_xx_flush_fe            (rtu_yy_xx_flush_fe           ),
  .vidu_rtu_no_op                (vidu_rtu_no_op               ),
  .vlsu_rtu_vl_updt_data         (vlsu_rtu_vl_updt_data        ),
  .vlsu_rtu_vl_updt_vld          (vlsu_rtu_vl_updt_vld         ),
  .vpu_rtu_ex1_cmplt             (vpu_rtu_ex1_cmplt            ),
  .vpu_rtu_ex1_cmplt_dp          (vpu_rtu_ex1_cmplt_dp         ),
  .vpu_rtu_ex1_fp_dirty          (vpu_rtu_ex1_fp_dirty         ),
  .vpu_rtu_ex1_vec_dirty         (vpu_rtu_ex1_vec_dirty        ),
  .vpu_rtu_fflag                 (vpu_rtu_fflag                ),
  .vpu_rtu_fflag_vld             (vpu_rtu_fflag_vld            ),
  .vpu_rtu_gpr_wb_data           (vpu_rtu_gpr_wb_data          ),
  .vpu_rtu_gpr_wb_index          (vpu_rtu_gpr_wb_index         ),
  .vpu_rtu_gpr_wb_req            (vpu_rtu_gpr_wb_req           ),
  .vpu_rtu_no_op                 (vpu_rtu_no_op                )
);

endmodule
